module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, StoB_REQ4_n, StoB_REQ5_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoS_ACK4_n, BtoS_ACK5_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, SLC2_n, jx0_n, jx1_n, jx2_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844f9d;
  wire v856422;
  wire v854b7c;
  wire v855fdf;
  wire v8a32ba;
  wire v856710;
  wire v857785;
  wire v8a3097;
  wire v857866;
  wire v85531b;
  wire v8a3151;
  wire v844f9f;
  wire v8a2972;
  wire v876d51;
  wire v854b1e;
  wire v857a31;
  wire v8a336c;
  wire v883730;
  wire v8a2d62;
  wire v854b2f;
  wire v85635c;
  wire v8a331b;
  wire v8575b3;
  wire v86f89c;
  wire v85523e;
  wire v855c3e;
  wire v856c80;
  wire v85628e;
  wire v8a3023;
  wire v857421;
  wire v8a31b7;
  wire v855748;
  wire v8a3260;
  wire v854a11;
  wire v8a308c;
  wire v8a2935;
  wire v8a3140;
  wire v8558ad;
  wire v854ffe;
  wire v8617fe;
  wire v8a3176;
  wire v8a3052;
  wire v844f9b;
  wire v88ab81;
  wire v8a3032;
  wire v8a30f6;
  wire v855ef6;
  wire v8558fe;
  wire v85778e;
  wire v8a31ca;
  wire v8a29d7;
  wire v8a3334;
  wire v8a30b8;
  wire v8a29eb;
  wire v8a3322;
  wire v856799;
  wire v8558e6;
  wire v844f99;
  wire v856c06;
  wire v8555ef;
  wire v857619;
  wire v855d5e;
  wire v8a3226;
  wire v8a31c5;
  wire v855865;
  wire v844f97;
  wire v8a30b3;
  wire v8a30b4;
  wire v8a33da;
  wire v86624f;
  wire v8555a0;
  wire v8a31c7;
  wire v8568be;
  wire v85a4b3;
  wire v85745e;
  wire v8a2a7f;
  wire v87116b;
  wire v85576e;
  wire v8a31e2;
  wire v857a21;
  wire v854138;
  wire v8579cf;
  wire v856111;
  wire v8550f3;
  wire v854b71;
  wire v8a32ea;
  wire v856863;
  wire v8a3282;
  wire v8a3042;
  wire v8679b5;
  wire v856e26;
  wire v8a33cd;
  wire v8a2489;
  wire v868cba;
  wire v896275;
  wire v855df9;
  wire v8a305b;
  wire v8a3286;
  wire v8960f3;
  wire v8a28b9;
  wire v8a2e89;
  wire v8a33c7;
  wire v87d011;
  wire v8552de;
  wire v8a312b;
  wire v855cb6;
  wire v87119a;
  wire v855501;
  wire v8a2d0e;
  wire v87734d;
  wire v8a30c4;
  wire v854b24;
  wire v854b5f;
  wire v85614f;
  wire v8a30e9;
  wire v855221;
  wire v856b4c;
  wire v8a3339;
  wire v8a32e8;
  wire v8a296b;
  wire v855d70;
  wire v86a9e8;
  wire v8a331a;
  wire v8a288c;
  wire v8a2c6b;
  wire v888ecd;
  wire v8557be;
  wire v8559ce;
  wire v854edc;
  wire v8a33de;
  wire v85510d;
  wire v85ecbc;
  wire v867ef3;
  wire v85eb80;
  wire v8a333c;
  wire v8a32eb;
  wire v85634e;
  wire v8a3272;
  wire v8557a6;
  wire v8a323a;
  wire v8a2b42;
  wire v85577c;
  wire v8a31ab;
  wire v859301;
  wire v8573d3;
  wire v855386;
  wire v855658;
  wire v8558d2;
  wire v8a300d;
  wire v8a30c1;
  wire v8a33c0;
  wire v85743a;
  wire v8a29cd;
  wire v8a3154;
  wire v8a308f;
  wire v8a33b0;
  wire v8a3026;
  wire v85504a;
  wire v8a3062;
  wire v8a3117;
  wire v856653;
  wire v856903;
  wire v85ecec;
  wire v871154;
  wire v8703da;
  wire v8a30d1;
  wire v85640f;
  wire v8a3088;
  wire v8557cd;
  wire v8a2b29;
  wire v8a3171;
  wire v857a8c;
  wire v88abc1;
  wire v8a32d8;
  wire v8558ef;
  wire v8a321c;
  wire v8a3075;
  wire v8a3179;
  wire v87532a;
  wire v8a30b7;
  wire v8575a5;
  wire v8553d5;
  wire v8a3182;
  wire v86aa3d;
  wire v89614f;
  wire v854c39;
  wire v8564e4;
  wire v85ab2f;
  wire v8565ef;
  wire v8a3346;
  wire v8a33e5;
  wire v8557f8;
  wire v855af2;
  wire v8a3187;
  wire v8a3236;
  wire v8711bb;
  wire v8a3302;
  wire v85554e;
  wire v855957;
  wire v8a308b;
  wire v8961d4;
  wire v844fad;
  wire v855f5b;
  wire v85741f;
  wire v8a3089;
  wire v8a31c8;
  wire v87c759;
  wire v85e22c;
  wire v8a2fba;
  wire v8685f8;
  wire v856d89;
  wire v8a29a5;
  wire v8a3265;
  wire v854ff9;
  wire v8a33d9;
  wire v854b6c;
  wire v8558ec;
  wire v855eb2;
  wire v8a315d;
  wire v854e55;
  wire v8a30fe;
  wire v8a327d;
  wire v8a3327;
  wire v8a2a54;
  wire v85aaf7;
  wire v8a332e;
  wire v8a29c6;
  wire v85528e;
  wire v8a31a7;
  wire v8562b9;
  wire v855d7a;
  wire v855d2c;
  wire v855b2d;
  wire v8a29f8;
  wire v8a30ef;
  wire v8558fa;
  wire v8563ed;
  wire v8a289a;
  wire v85570e;
  wire v854ee4;
  wire v8a24df;
  wire v8a283f;
  wire v8a3147;
  wire v856c7e;
  wire v86da55;
  wire v861d68;
  wire v857932;
  wire v8552c8;
  wire v855065;
  wire v8562af;
  wire v856441;
  wire v855492;
  wire v86917e;
  wire v8565de;
  wire v871138;
  wire v8a3183;
  wire v8579da;
  wire v8a310e;
  wire v8a2ef0;
  wire v854a55;
  wire v8a3066;
  wire v854f1c;
  wire v856543;
  wire v854e7c;
  wire v8a2bf7;
  wire v8a2ffa;
  wire v856417;
  wire v89626e;
  wire v855d34;
  wire v8a31ac;
  wire v8579fd;
  wire v85594d;
  wire v8a3275;
  wire v85694d;
  wire v8a3300;
  wire v8565b9;
  wire v855ed8;
  wire v8a314d;
  wire v856781;
  wire v856374;
  wire v8565a7;
  wire v854f04;
  wire v856e4a;
  wire v8a329d;
  wire v8a2dfb;
  wire v857583;
  wire v8579f4;
  wire v855e0d;
  wire v85756f;
  wire v856535;
  wire v8a3415;
  wire v856195;
  wire v8561a3;
  wire v855786;
  wire v854a35;
  wire v854d07;
  wire v855bec;
  wire v855b6e;
  wire v856b86;
  wire v855505;
  wire v85768c;
  wire v854ccd;
  wire v8575fe;
  wire v875b8c;
  wire v8560a3;
  wire v8a31c0;
  wire v86179a;
  wire v85682b;
  wire v855a8a;
  wire v8a312e;
  wire v855033;
  wire v8a3227;
  wire v8a3120;
  wire v856b6b;
  wire v8a3143;
  wire v8550e8;
  wire v85607f;
  wire v8a3108;
  wire v85aac2;
  wire v8a2837;
  wire v854d1f;
  wire v8836e5;
  wire v8a291b;
  wire v896167;
  wire v861800;
  wire v883cae;
  wire v856e02;
  wire v8a2f1e;
  wire v8573f3;
  wire v88abca;
  wire v8a3342;
  wire v8575aa;
  wire v8a30e1;
  wire v855845;
  wire v8553df;
  wire v85a3c4;
  wire v8a33bc;
  wire v856ab0;
  wire v855fec;
  wire v8a305e;
  wire v8a0e69;
  wire v844fa1;
  wire v844fa0;
  wire v855b05;
  wire v856562;
  wire v856af3;
  wire v871675;
  wire v852505;
  wire v8563c1;
  wire v8a334f;
  wire v88372d;
  wire v8962e0;
  wire v8a30c9;
  wire v8961ac;
  wire v844f95;
  wire v8a2fd5;
  wire v8a284d;
  wire v8a317f;
  wire v8a329f;
  wire v8a3329;
  wire v86f537;
  wire v8a3211;
  wire v85ed68;
  wire v883725;
  wire v8a332c;
  wire v89624b;
  wire v8a3058;
  wire v856992;
  wire v8a33be;
  wire v857a0d;
  wire v85eda6;
  wire v8a3132;
  wire v88ab87;
  wire v8a3045;
  wire v86aa63;
  wire v855db1;
  wire v8a3107;
  wire v8a2a91;
  wire v855acd;
  wire v85778c;
  wire v8a3142;
  wire v8a326c;
  wire v8a33c1;
  wire v86c421;
  wire v856ab3;
  wire v855e00;
  wire v8a3081;
  wire v857692;
  wire v8a2cab;
  wire v8576bc;
  wire v8a294c;
  wire v86c9ca;
  wire v883cb2;
  wire v85544e;
  wire v8559ee;
  wire v8a2e46;
  wire v860093;
  wire v85699f;
  wire v86a9cb;
  wire v8a3235;
  wire v8a311d;
  wire v8a3317;
  wire v856aac;
  wire v855426;
  wire v8a30e7;
  wire v8a334a;
  wire v8a2d94;
  wire v88375a;
  wire v89625f;
  wire v8a3318;
  wire v88b742;
  wire v896107;
  wire v85a3a7;
  wire v8a328b;
  wire v85613d;
  wire v856cd1;
  wire v8a297d;
  wire v8a307a;
  wire v8a2c65;
  wire v8556ec;
  wire v857b51;
  wire v844fc1;
  wire v8a2d10;
  wire v8549e6;
  wire v873280;
  wire v86cbc9;
  wire v854fc1;
  wire v85743c;
  wire v855998;
  wire v873756;
  wire v8a2fa9;
  wire v855bf8;
  wire v8a3367;
  wire v8962ff;
  wire v844fbd;
  wire v844fbf;
  wire v855db2;
  wire v8a30f8;
  wire v8a30dc;
  wire v8a28a9;
  wire v8a32e1;
  wire v8a32ef;
  wire v8a3320;
  wire v88ea49;
  wire v8a3043;
  wire v8a2eb6;
  wire v85610f;
  wire v85540d;
  wire v8a2a8c;
  wire v8a2f7a;
  wire v8a311e;
  wire v8559f8;
  wire v89fcfa;
  wire v858bbc;
  wire v8a30cf;
  wire v87bbfb;
  wire v856648;
  wire v8a3163;
  wire v857b70;
  wire v856982;
  wire v857624;
  wire v876345;
  wire v854fc7;
  wire v8a3027;
  wire v856c9f;
  wire v88373a;
  wire v8a330f;
  wire v883733;
  wire v8a306b;
  wire v8961a6;
  wire v856730;
  wire v857595;
  wire v8a3167;
  wire v8a32bd;
  wire v896294;
  wire v8a31e3;
  wire v8549ca;
  wire v85618d;
  wire v856c72;
  wire v854b14;
  wire v856abb;
  wire v8a33a5;
  wire v854fcb;
  wire v8556a7;
  wire v856c11;
  wire v888edb;
  wire v855311;
  wire v8a32f4;
  wire v8a3350;
  wire v8551d0;
  wire v86f804;
  wire v855cd0;
  wire v8a338c;
  wire v85606a;
  wire v8a3086;
  wire v8711c0;
  wire v855c79;
  wire v85532e;
  wire v8a322d;
  wire v8961a8;
  wire v8711d9;
  wire v872af1;
  wire v8a3128;
  wire v85ed30;
  wire v8a334e;
  wire v857aed;
  wire v86938f;
  wire v854feb;
  wire v85ed6f;
  wire v8711cf;
  wire v8a3377;
  wire v8a2b0e;
  wire v854ed3;
  wire v8a3096;
  wire v8a31b9;
  wire v883709;
  wire v8a336a;
  wire v88abed;
  wire v8a31ba;
  wire v856ac3;
  wire v8a2c94;
  wire v856438;
  wire v8a3112;
  wire v8573b7;
  wire v8a32a7;
  wire v8a3144;
  wire v8a3099;
  wire v8557b8;
  wire v85ab66;
  wire v8a33d5;
  wire v855268;
  wire v85765d;
  wire v8574eb;
  wire v855361;
  wire v86c425;
  wire v8560c5;
  wire v856651;
  wire v856786;
  wire v8567c7;
  wire v8a3354;
  wire v8a314b;
  wire v8a331c;
  wire v855735;
  wire v8a2d1f;
  wire v856670;
  wire v8a32a4;
  wire v854ae3;
  wire v8a321d;
  wire v857547;
  wire v89612f;
  wire v856467;
  wire v8a32fd;
  wire v856e00;
  wire v857880;
  wire v873869;
  wire v8a3074;
  wire v8a3340;
  wire v8a31b3;
  wire v8a3158;
  wire v8a3152;
  wire v856cee;
  wire v8a30bf;
  wire v857694;
  wire v85601f;
  wire v85524b;
  wire v855681;
  wire v8565ba;
  wire v854188;
  wire v8552f8;
  wire v8a30ac;
  wire v856df1;
  wire v8a3307;
  wire v8a31b1;
  wire v85edf0;
  wire v8a299a;
  wire v856c23;
  wire v854ae5;
  wire v876a61;
  wire v855879;
  wire v8550be;
  wire v8836fc;
  wire v8560bc;
  wire v857651;
  wire v8a3355;
  wire v8a3330;
  wire v8a2dc2;
  wire v8a3249;
  wire v8a331e;
  wire v8a30ce;
  wire v86a9cf;
  wire v8a338e;
  wire v855e36;
  wire v855f60;
  wire v8a318e;
  wire v8a2893;
  wire v85687a;
  wire v8a313d;
  wire v855791;
  wire v8557e6;
  wire v854ef2;
  wire v8553de;
  wire v856102;
  wire v856761;
  wire v855418;
  wire v854d3e;
  wire v8a33c4;
  wire v85759c;
  wire v8556cb;
  wire v857689;
  wire v855c38;
  wire v867273;
  wire v8a2b16;
  wire v8a3184;
  wire v85754a;
  wire v8560c6;
  wire v857a0c;
  wire v855c3a;
  wire v8573e8;
  wire v8a3242;
  wire v8a323e;
  wire v85586d;
  wire v8a3193;
  wire v8a32a9;
  wire v8a32af;
  wire v857b42;
  wire v8a320d;
  wire v85509f;
  wire v8a317b;
  wire v8a2bd1;
  wire v86a9c5;
  wire v8a31d5;
  wire v856047;
  wire v87c729;
  wire v8532c4;
  wire v868e49;
  wire v856636;
  wire v855078;
  wire v8567b5;
  wire v8a3229;
  wire v85663b;
  wire v856b2a;
  wire v8a31cc;
  wire v8a311b;
  wire v8551a3;
  wire v8a2ce0;
  wire v855c86;
  wire v896248;
  wire v8a32cc;
  wire v854ba4;
  wire v8a338b;
  wire v855bae;
  wire v8a3156;
  wire v8a3387;
  wire v85646a;
  wire v85793b;
  wire v857418;
  wire v88ab43;
  wire v8a3214;
  wire v85ed1a;
  wire v8a2bb0;
  wire v8a3038;
  wire v8a30ba;
  wire v8a2c17;
  wire v86178d;
  wire v856443;
  wire v85660e;
  wire v8a2fd8;
  wire v8541e8;
  wire v85762e;
  wire v8a2ee2;
  wire v865746;
  wire v8a313e;
  wire v8a3185;
  wire v856d80;
  wire v8574ee;
  wire v855631;
  wire v8558ea;
  wire v8578b4;
  wire v85690e;
  wire v8a30be;
  wire v855850;
  wire v855182;
  wire v8a32e2;
  wire v8a322c;
  wire v8a310d;
  wire v856784;
  wire v8a287f;
  wire v8a3299;
  wire v877887;
  wire v8a339d;
  wire v88a46b;
  wire v8617be;
  wire v8554bf;
  wire v8a3325;
  wire v855bdb;
  wire v8a303b;
  wire v855564;
  wire v85ab2a;
  wire v8a306e;
  wire v8a3301;
  wire v856431;
  wire v8a3206;
  wire v854c99;
  wire v8a2c75;
  wire v8a31ae;
  wire v8a3049;
  wire v8551ba;
  wire v8a3251;
  wire v8a3245;
  wire v8a30b0;
  wire v8a3160;
  wire v856723;
  wire v8a3364;
  wire v8a2fc5;
  wire v8561e1;
  wire v88a458;
  wire v8555b7;
  wire v856b1f;
  wire v8a3290;
  wire v855e40;
  wire v8a30bb;
  wire v8a31dc;
  wire v85548d;
  wire v8556fc;
  wire v8563d8;
  wire v876637;
  wire v855700;
  wire v856144;
  wire v856991;
  wire v8a328e;
  wire v8a33d3;
  wire v8a3363;
  wire v8a2f07;
  wire v8a30c2;
  wire v8a32cb;
  wire v8a2aed;
  wire v8a3101;
  wire v8a311c;
  wire v855cd9;
  wire v85677d;
  wire v8558cf;
  wire v8551dd;
  wire v8a29dc;
  wire v85586a;
  wire v8a3253;
  wire v8a32a3;
  wire v85d533;
  wire v856003;
  wire v857b78;
  wire v8562e3;
  wire v85eae9;
  wire v88ac2c;
  wire v8a32f8;
  wire v856af6;
  wire v854151;
  wire v8a3094;
  wire v8a3090;
  wire v871174;
  wire v8a303e;
  wire v8a304c;
  wire v8a31af;
  wire v8a0e17;
  wire v8a30b1;
  wire v85d4ae;
  wire v8a325f;
  wire v8a3380;
  wire v8a32ae;
  wire v8a3083;
  wire v854cf3;
  wire v854c4e;
  wire v855e1c;
  wire v8a33df;
  wire v8a2ff0;
  wire v855708;
  wire v8556c9;
  wire v8567ad;
  wire v857aee;
  wire v856a98;
  wire v8a3221;
  wire v8a30c3;
  wire v855d3a;
  wire v855c80;
  wire v854204;
  wire v855a47;
  wire v855283;
  wire v8a3022;
  wire v8a30dd;
  wire v8a30e0;
  wire v8a309d;
  wire v856256;
  wire v8a3321;
  wire v88a46f;
  wire v854aed;
  wire v8a2be7;
  wire v844fa3;
  wire v8a32fe;
  wire v85648f;
  wire v856945;
  wire v854f2f;
  wire v8a30ec;
  wire v86f7aa;
  wire v8550af;
  wire v883756;
  wire v856737;
  wire v883ce3;
  wire v844fa9;
  wire v8a3175;
  wire v8a30f7;
  wire v854e78;
  wire v8552ea;
  wire v856678;
  wire v8a31b8;
  wire v85bce8;
  wire v855d84;
  wire v8a3207;
  wire v8a32c0;
  wire v857a54;
  wire v8a2daf;
  wire v85be20;
  wire v854fd3;
  wire v8566c4;
  wire v854cc4;
  wire v8a0dfa;
  wire v8a3002;
  wire v8a282b;
  wire v855a2a;
  wire v8a30a5;
  wire v8a302e;
  wire v8a3035;
  wire v8738de;
  wire v856bea;
  wire v8a3273;
  wire v88abf3;
  wire v856545;
  wire v855edf;
  wire v8a3258;
  wire v8a315b;
  wire v8960fd;
  wire v856926;
  wire v8711ac;
  wire v8566b8;
  wire v856828;
  wire v876d41;
  wire v8567aa;
  wire v8662d9;
  wire v855aec;
  wire v856966;
  wire v85aae3;
  wire v856434;
  wire v8a333b;
  wire v8a33ae;
  wire v86a9f3;
  wire v8a3196;
  wire v8558f4;
  wire v88a469;
  wire v8a3284;
  wire v856e3f;
  wire v8a3244;
  wire v8a32c6;
  wire v8617f7;
  wire v8a310a;
  wire v855d7f;
  wire v85786a;
  wire v85e7e0;
  wire v8a309b;
  wire v8a335a;
  wire v85a4b2;
  wire v858911;
  wire v854aa0;
  wire v856d91;
  wire v855f55;
  wire v8a2486;
  wire v8558cb;
  wire v8a3388;
  wire v85665d;
  wire v85528a;
  wire v8a2c6e;
  wire v86dd6d;
  wire v8a3040;
  wire v8a28d0;
  wire v8a2d12;
  wire v85579f;
  wire v8a3016;
  wire v88ab99;
  wire v8a312d;
  wire v86a9eb;
  wire v8556d0;
  wire v8a3305;
  wire v8a3345;
  wire v855870;
  wire v8a3091;
  wire v855de8;
  wire v8a3079;
  wire v8a3110;
  wire v8a24b8;
  wire v855ebf;
  wire v85566d;
  wire v8a2bb4;
  wire v8a30cd;
  wire v8a320e;
  wire v8a2e76;
  wire v855e45;
  wire v8556bc;
  wire v8a32da;
  wire v866b88;
  wire v855a61;
  wire v8a32d0;
  wire v85edc8;
  wire v854a23;
  wire v8a28de;
  wire v8a0de5;
  wire v855a4d;
  wire v856db6;
  wire v883775;
  wire v8560ea;
  wire v8a3082;
  wire v8a3314;
  wire v8573cd;
  wire v85413e;
  wire v8a337f;
  wire v856883;
  wire v8541c6;
  wire v85ab2e;
  wire v854a89;
  wire v854a17;
  wire v8561e7;
  wire v856b69;
  wire v8567ec;
  wire v8a3170;
  wire v844fe7;
  wire v854d33;
  wire v8a3166;
  wire v8a3135;
  wire v88abdb;
  wire v855ffb;
  wire v8a2b82;
  wire v8a30eb;
  wire v86aa28;
  wire v8a30d8;
  wire v8541a9;
  wire v856026;
  wire v8a3332;
  wire v883cad;
  wire v8a31d2;
  wire v8a32df;
  wire v856262;
  wire v855c9e;
  wire v85676f;
  wire v8a315e;
  wire v89fce5;
  wire v85575f;
  wire v870d30;
  wire v857783;
  wire v856253;
  wire v8a2dfa;
  wire v86eb76;
  wire v856b26;
  wire v8a335b;
  wire v85ec27;
  wire v8a2b44;
  wire v855e0c;
  wire v856432;
  wire v88abd1;
  wire v857a7a;
  wire v844fb1;
  wire v856302;
  wire v8a2d78;
  wire v8a33ce;
  wire v86aa4d;
  wire v8a3033;
  wire v8a309a;
  wire v8552b8;
  wire v85617a;
  wire v8a2dbf;
  wire v856041;
  wire v8a33b3;
  wire v8a319c;
  wire v869f3f;
  wire v855e0e;
  wire v8a3208;
  wire v8a30b6;
  wire v8573a4;
  wire v8a31f4;
  wire v86b41a;
  wire v8a0e03;
  wire v855a7a;
  wire v854b1a;
  wire v883710;
  wire v8a30fd;
  wire v856e34;
  wire v8579a9;
  wire v856e7b;
  wire v855014;
  wire v8a3159;
  wire v8566e6;
  wire v854c44;
  wire v8a337e;
  wire v857af8;
  wire v8a2f6b;
  wire v856007;
  wire v8a3194;
  wire v855016;
  wire v8550a0;
  wire v8a328d;
  wire v8a3031;
  wire v854cad;
  wire v8a3181;
  wire v87c763;
  wire v8565c6;
  wire v857649;
  wire v8a2d89;
  wire v8a3189;
  wire v8a2824;
  wire v883c9a;
  wire v8a2e8b;
  wire v867269;
  wire v856c36;
  wire v88ac3b;
  wire v8a2898;
  wire v85aab4;
  wire v8a3233;
  wire v8557e1;
  wire v8a33aa;
  wire v8a30a3;
  wire v85651f;
  wire v85797a;
  wire v8a327e;
  wire v8a319e;
  wire v8a30ab;
  wire v8564e9;
  wire v8550c7;
  wire v856130;
  wire v857b8b;
  wire v8a3219;
  wire v8a326d;
  wire v8a302f;
  wire v883759;
  wire v8a33b2;
  wire v8a2485;
  wire v856352;
  wire v85644e;
  wire v855185;
  wire v8a33cf;
  wire v8a3262;
  wire v855dee;
  wire v855c77;
  wire v8a30f0;
  wire v8554e5;
  wire v8a302d;
  wire v855b1d;
  wire v857a4d;
  wire v8568ac;
  wire v883cb8;
  wire v8a30b5;
  wire v857775;
  wire v854f98;
  wire v8a30af;
  wire v8a3234;
  wire v8554d7;
  wire v8a30fb;
  wire v8a304b;
  wire v8a30aa;
  wire v8a307b;
  wire v85623b;
  wire v8a2b13;
  wire v855218;
  wire v8a2ef9;
  wire v857aaa;
  wire v855ac2;
  wire v88abaa;
  wire v8574ef;
  wire v855565;
  wire v8a30e6;
  wire v8559e7;
  wire v8a30a6;
  wire v855fac;
  wire v8a33b1;
  wire v8a3198;
  wire v86aa1f;
  wire v85562c;
  wire v85a3a3;
  wire v855e5a;
  wire v857a65;
  wire v8a3223;
  wire v85e12c;
  wire v87c76f;
  wire v844fab;
  wire v856553;
  wire v8552e8;
  wire v85698e;
  wire v855e66;
  wire v8a336d;
  wire v86aa4b;
  wire v8a33c2;
  wire v8a3077;
  wire v85698c;
  wire v8a316d;
  wire v86aa49;
  wire v8a3285;
  wire v8579f3;
  wire v88b745;
  wire v8a333a;
  wire v8564d2;
  wire v8a3241;
  wire v8a3292;
  wire v8a2d93;
  wire v856bc0;
  wire v8a3178;
  wire v855397;
  wire v8a3361;
  wire v8a3392;
  wire v8a3263;
  wire v8a3129;
  wire v8a2c6c;
  wire v8a2d29;
  wire v857ad0;
  wire v8a3098;
  wire v855c08;
  wire v8a3386;
  wire v8552ac;
  wire v85795e;
  wire v8a0de9;
  wire v8a3313;
  wire v854be5;
  wire v855196;
  wire v86007c;
  wire v8554b2;
  wire v855f7c;
  wire v855a02;
  wire v8a332a;
  wire v8555d3;
  wire v855583;
  wire v8a31cd;
  wire v88a44b;
  wire v8a2e94;
  wire v855533;
  wire v896162;
  wire v8550a1;
  wire v856be3;
  wire v8a302a;
  wire v8a32c4;
  wire v856ad7;
  wire v8738b2;
  wire v8a3362;
  wire v854fa7;
  wire v8579c7;
  wire v860488;
  wire v8a29e3;
  wire v877670;
  wire v896106;
  wire v85413d;
  wire v85499f;
  wire v856023;
  wire v856d52;
  wire v8a338f;
  wire v896289;
  wire v8a329c;
  wire v855fb5;
  wire v88abc5;
  wire v855c02;
  wire v8a321f;
  wire v855f43;
  wire v8a30de;
  wire v8a30b2;
  wire v8576d5;
  wire v8a304e;
  wire v8a2fb0;
  wire v8a2e00;
  wire v856731;
  wire v89629f;
  wire v8a2958;
  wire v8a3053;
  wire v8557f6;
  wire v8a2d8d;
  wire v8a31d1;
  wire v856801;
  wire v8a3389;
  wire v856c01;
  wire v8a328a;
  wire v8a2a74;
  wire v854f8b;
  wire v857979;
  wire v855a09;
  wire v8a31ad;
  wire v855b2c;
  wire v8a2cc7;
  wire v8541e6;
  wire v8a3347;
  wire v8574e2;
  wire v855060;
  wire v85659e;
  wire v85658a;
  wire v855002;
  wire v8a31aa;
  wire v854cb1;
  wire v8a31d0;
  wire v8a2a85;
  wire v8a295f;
  wire v8a31bb;
  wire v8a30fc;
  wire v8a0e3c;
  wire v8566b6;
  wire v8a3294;
  wire v8a315c;
  wire v855cc1;
  wire v8a30d5;
  wire v855ab2;
  wire v854d31;
  wire v855b5d;
  wire v855f89;
  wire v855d3e;
  wire v8a3080;
  wire v888ec4;
  wire v8a3287;
  wire v8a32a1;
  wire v8a287d;
  wire v8a2e77;
  wire v856197;
  wire v8562f8;
  wire v8a320a;
  wire v855ebc;
  wire v8a2c53;
  wire v855d44;
  wire v8962f6;
  wire v857414;
  wire v8a31e6;
  wire v8a31c6;
  wire v8a3118;
  wire v855c15;
  wire v856b13;
  wire v8a2fce;
  wire v8554f7;
  wire v855ddf;
  wire v8a317d;
  wire v855fb0;
  wire v85ab14;
  wire v88abc3;
  wire v854a07;
  wire v8a3131;
  wire v85500c;
  wire v8a2c62;
  wire v856c8d;
  wire v85554c;
  wire v85edf1;
  wire v85509b;
  wire v873fa6;
  wire v8a2f46;
  wire v855254;
  wire v857969;
  wire v857534;
  wire v855c6b;
  wire v855eb3;
  wire v856624;
  wire v8a3315;
  wire v871051;
  wire v854c82;
  wire v8a2b19;
  wire v85555c;
  wire v8552b4;
  wire v8962c7;
  wire v8a2ae0;
  wire v867265;
  wire v8a30e5;
  wire v855780;
  wire v8551f8;
  wire v854fff;
  wire v8a3270;
  wire v8a332b;
  wire v8a33d8;
  wire v855faf;
  wire v855ba9;
  wire v854a0a;
  wire v87116a;
  wire v854a53;
  wire v8a337d;
  wire v8a320f;
  wire v8a306f;
  wire v855df1;
  wire v8559aa;
  wire v855d45;
  wire v85543e;
  wire v855398;
  wire v856270;
  wire v85576d;
  wire v8a31a8;
  wire v85565b;
  wire v8a2e72;
  wire v855653;
  wire v855858;
  wire v8a3372;
  wire v854a06;
  wire v86fe32;
  wire v8551f9;
  wire v856063;
  wire v8a3279;
  wire v856e74;
  wire v855ee6;
  wire v854f97;
  wire v857917;
  wire v870eba;
  wire v8a339a;
  wire v8a30bd;
  wire v8560aa;
  wire v8a3164;
  wire v85796e;
  wire v856835;
  wire v855298;
  wire v8a31b6;
  wire v8a3336;
  wire v8a30c5;
  wire v855d6a;
  wire v8a2448;
  wire v857543;
  wire v8a2b63;
  wire v8a32d3;
  wire v87d033;
  wire v855e79;
  wire v8560fa;
  wire v8a324c;
  wire v873613;
  wire v8a3376;
  wire v855941;
  wire v8a2ec1;
  wire v856e47;
  wire v8a31f2;
  wire v8a32ce;
  wire v8a28c6;
  wire v8a329e;
  wire v870ea7;
  wire v8a331f;
  wire v8a33c6;
  wire v8a31ee;
  wire v85508c;
  wire v85683b;
  wire v8a336e;
  wire v85ab44;
  wire v8a0e4e;
  wire v85d977;
  wire v856cce;
  wire v8617d4;
  wire v856b8f;
  wire v8961a7;
  wire v854fe3;
  wire v873853;
  wire v855f3f;
  wire v8a3326;
  wire v856dec;
  wire v855069;
  wire v8a31a1;
  wire v8a3358;
  wire v8566ad;
  wire v8a3225;
  wire v854cbb;
  wire v854b8e;
  wire v8a327a;
  wire v8556c1;
  wire v855709;
  wire v857487;
  wire v8a3197;
  wire v8a31a9;
  wire v8a309e;
  wire v855ce1;
  wire v856b58;
  wire v856884;
  wire v855414;
  wire v8a3149;
  wire v87c747;
  wire v896174;
  wire v8a3106;
  wire v8a31a2;
  wire v854b5e;
  wire v856901;
  wire v8a32fb;
  wire v8559bc;
  wire v8a28af;
  wire v855ea7;
  wire v8a3228;
  wire v87116e;
  wire v856bfd;
  wire v856264;
  wire v86aa64;
  wire v8a3232;
  wire v854bcd;
  wire v854b33;
  wire v8a29ad;
  wire v856288;
  wire v87c743;
  wire v855bc8;
  wire v85a071;
  wire v855046;
  wire v8a324a;
  wire v8a2f21;
  wire v869886;
  wire v854c76;
  wire v856790;
  wire v87d020;
  wire v85751a;
  wire v85581e;
  wire v8569e1;
  wire v854c5c;
  wire v861784;
  wire v8568b1;
  wire v856075;
  wire v85522d;
  wire v8a3289;
  wire v8a31bd;
  wire v8a247a;
  wire v85621e;
  wire v8a3360;
  wire v8a3050;
  wire v88abb8;
  wire v8a31fa;
  wire v855783;
  wire v85eb9f;
  wire v85edeb;
  wire v857b65;
  wire v8a3393;
  wire v8a0e4f;
  wire v870eb8;
  wire v8961ce;
  wire v855001;
  wire v8a2d44;
  wire v8569fe;
  wire v8573ee;
  wire v854f52;
  wire v85791e;
  wire v8a3130;
  wire v8553e6;
  wire v873899;
  wire v85be78;
  wire v857b07;
  wire v85aad7;
  wire v8551c8;
  wire v856b54;
  wire v854f90;
  wire v854c5b;
  wire v8a31ed;
  wire v8558d9;
  wire v8553cf;
  wire v8a24a6;
  wire v8a2d5b;
  wire v8a329b;
  wire v856176;
  wire v8a31e4;
  wire v8a31b2;
  wire v89cb27;
  wire v856556;
  wire v8a30e2;
  wire v8a30d3;
  wire v855f95;
  wire v8a3250;
  wire v8a3153;
  wire v8654fb;
  wire v8a3030;
  wire v8a330a;
  wire v85678b;
  wire v854fe9;
  wire v8a3036;
  wire v856639;
  wire v8a3379;
  wire v854e79;
  wire v8560f5;
  wire v857452;
  wire v8a3395;
  wire v856a09;
  wire v8558a0;
  wire v855a9b;
  wire v85edc7;
  wire v8a304f;
  wire v8a2e4a;
  wire v856e5f;
  wire v855c5f;
  wire v8567b8;
  wire v855912;
  wire v8a336b;
  wire v855d52;
  wire v854e8e;
  wire v8a313f;
  wire v856acb;
  wire v8630d3;
  wire v855600;
  wire v857731;
  wire v855790;
  wire v8a31c1;
  wire v856062;
  wire v89caa5;
  wire v855531;
  wire v856bdb;
  wire v8a31f3;
  wire v88ab9d;
  wire v857469;
  wire v8a32a6;
  wire v8a3338;
  wire v8554aa;
  wire v8552f4;
  wire v863beb;
  wire v8a31d8;
  wire v8a3309;
  wire v8a32b6;
  wire v8a3391;
  wire v85509e;
  wire v8a31ea;
  wire v854a8f;
  wire v8a2ddc;
  wire v8566d2;
  wire v85a48b;
  wire v85ecc8;
  wire v88ab6c;
  wire v8a329a;
  wire v8a2c28;
  wire v8549ee;
  wire v855b24;
  wire v8a3239;
  wire v8569b3;
  wire v8a2cce;
  wire v855acb;
  wire v8a323b;
  wire v8a3288;
  wire v854bf7;
  wire v856e2b;
  wire v8549db;
  wire v8774cb;
  wire v854a71;
  wire v8560ec;
  wire v8a3269;
  wire v8a339b;
  wire v8a33ec;
  wire v854eb2;
  wire v8a2fe8;
  wire v856c4f;
  wire v856df4;
  wire v856575;
  wire v8a32b8;
  wire v855e06;
  wire v8a3303;
  wire v855114;
  wire v8564c9;
  wire v856e10;
  wire v856e0b;
  wire v8738ae;
  wire v8a3220;
  wire v8a2e42;
  wire v85605e;
  wire v87c300;
  wire v855314;
  wire v85a137;
  wire v8a31e5;
  wire v8a24c7;
  wire v8a243e;
  wire v857521;
  wire v8a0e55;
  wire v8a3203;
  wire v856313;
  wire v855147;
  wire v8549e9;
  wire v8a32b3;
  wire v8560ff;
  wire v856847;
  wire v854ed7;
  wire v883754;
  wire v855e27;
  wire v8a2f17;
  wire v8a3044;
  wire v8576c3;
  wire v8a333f;
  wire v8549c4;
  wire v855126;
  wire v8961cb;
  wire v855894;
  wire v854d20;
  wire v870ea9;
  wire v8566e1;
  wire v8a31b0;
  wire v85746e;
  wire v8a31fb;
  wire v888ed9;
  wire v85419c;
  wire v855674;
  wire v8549fe;
  wire v8551da;
  wire v8960ee;
  wire v85749f;
  wire v8711df;
  wire v8a2fac;
  wire v8567a3;
  wire v8a3150;
  wire v8a326b;
  wire v856c57;
  wire v8553e7;
  wire v8559d2;
  wire v8a2a3d;
  wire v865fb9;
  wire v854edf;
  wire v8a3116;
  wire v86c364;
  wire v8a3237;
  wire v855739;
  wire v856497;
  wire v876d53;
  wire v8a2bfd;
  wire v88371a;
  wire v8a3243;
  wire v8541c3;
  wire v856aa1;
  wire v8a3217;
  wire v8a2e9b;
  wire v8a3115;
  wire v8a0e0a;
  wire v8a318a;
  wire v856436;
  wire v8a32b9;
  wire v8a3278;
  wire v8a3210;
  wire v854b17;
  wire v8a2cbd;
  wire v8a2e43;
  wire v883741;
  wire v8a33db;
  wire v8a3222;
  wire v856489;
  wire v854994;
  wire v8a31bc;
  wire v857727;
  wire v85747f;
  wire v854d01;
  wire v87e83a;
  wire v8a33ac;
  wire v88ab84;
  wire v8a304d;
  wire v8a3095;
  wire v8a3202;
  wire v8a3398;
  wire v8575b5;
  wire v855ae0;
  wire v8a2891;
  wire v854988;
  wire v8568b8;
  wire v85531c;
  wire v87c6f7;
  wire v8574f8;
  wire v8a2f81;
  wire v8a32d7;
  wire v854b0e;
  wire v8a314c;
  wire v855d98;
  wire v8a325b;
  wire v855d54;
  wire v854a65;
  wire v856885;
  wire v8a283c;
  wire v854cd0;
  wire v85525c;
  wire v855e0f;
  wire v85555f;
  wire v854c40;
  wire v8a316b;
  wire v8a31ff;
  wire v8a2faa;
  wire v855a89;
  wire v88ab71;
  wire v8a2f9b;
  wire v8562a3;
  wire v856ad5;
  wire v8a3405;
  wire v8a3155;
  wire v8573a2;
  wire v856ad2;
  wire v8557b0;
  wire v8a3173;
  wire v8a307c;
  wire v8a31df;
  wire v8a31b5;
  wire v8550db;
  wire v8558d6;
  wire v8a3134;
  wire v855a66;
  wire v8a32d9;
  wire v878154;
  wire v8a24d1;
  wire v85be86;
  wire v8a2e1f;
  wire v866887;
  wire v844faf;
  wire v861796;
  wire v856705;
  wire v8574ba;
  wire v8a3186;
  wire v85681c;
  wire v855833;
  wire v855042;
  wire v8a31fe;
  wire v86e4e3;
  wire v8550b4;
  wire v854194;
  wire v87c725;
  wire v8a313a;
  wire v856871;
  wire v8a3025;
  wire v85522b;
  wire v855011;
  wire v8562d8;
  wire v856e7f;
  wire v8a3356;
  wire v854d35;
  wire v8a2da1;
  wire v8550fb;
  wire v85601a;
  wire v854f9b;
  wire v8a31dd;
  wire v8a326f;
  wire v8a30c7;
  wire v8a2c50;
  wire v8a2fa6;
  wire v85adee;
  wire v855edc;
  wire v855935;
  wire v87c707;
  wire v8a33e8;
  wire v857a91;
  wire v857a8e;
  wire v8a3268;
  wire v86b201;
  wire v854f20;
  wire v855ff1;
  wire v856bd6;
  wire v854eb5;
  wire v85520c;
  wire v8a33ad;
  wire v8a3200;
  wire v8a32c3;
  wire v8563cf;
  wire v8541c7;
  wire v855cfe;
  wire v8563a6;
  wire v856500;
  wire v855542;
  wire v8a3257;
  wire v85416e;
  wire v8a2a05;
  wire v85628f;
  wire v8549bd;
  wire v8a31d9;
  wire v855528;
  wire v8a330c;
  wire v8552c6;
  wire v8a3399;
  wire v8a3046;
  wire v8a315a;
  wire v85685d;
  wire v854eff;
  wire v8a3333;
  wire v855e7a;
  wire v85798c;
  wire v8a307d;
  wire v8a327f;
  wire v8a339f;
  wire v8a2479;
  wire v8a3070;
  wire v855b2b;
  wire v855fab;
  wire v8a2ff2;
  wire v855137;
  wire v857572;
  wire v8a3381;
  wire v8566bd;
  wire v8a3048;
  wire v8a2f08;
  wire v8962fa;
  wire v8a3397;
  wire v8a3267;
  wire v8560e2;
  wire v857674;
  wire v854ffa;
  wire v86a9dc;
  wire v856349;
  wire v8a3408;
  wire v883cb1;
  wire v8a32f2;
  wire v8578fc;
  wire v8a3246;
  wire v8a33af;
  wire v85675f;
  wire v8a3054;
  wire v8691ce;
  wire v855a8f;
  wire v8a2b95;
  wire v8a3261;
  wire v8a2bfa;
  wire v855ead;
  wire v855a6a;
  wire v856372;
  wire v86550e;
  wire v8a29d0;
  wire v8a321e;
  wire v8a2984;
  wire v85ab38;
  wire v856495;
  wire v8a2d5f;
  wire v8a3304;
  wire v855047;
  wire v8561c3;
  wire v86aa4a;
  wire v86e908;
  wire v8a31fd;
  wire v8a31f6;
  wire v8579f9;
  wire v8a302c;
  wire v8a2894;
  wire v85a4b4;
  wire v8a3293;
  wire v8617c9;
  wire v88ab9b;
  wire v873866;
  wire v8a31cb;
  wire v86d760;
  wire v85679c;
  wire v86180e;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg StoB_REQ4_p;
  input StoB_REQ4_n;
  reg StoB_REQ5_p;
  input StoB_REQ5_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoS_ACK4_p;
  output BtoS_ACK4_n;
  reg BtoS_ACK5_p;
  output BtoS_ACK5_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg SLC2_p;
  output SLC2_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  wire ENQ_n;
  wire SLC2_n;

assign v8a3338 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8a32a6;
assign v8a2d44 = jx2_p & v8a31fa | !jx2_p & !v855001;
assign v8a32da = jx2_p & v8556bc | !jx2_p & v844fa9;
assign v85aae3 = StoB_REQ0_p & v8a2b16 | !StoB_REQ0_p & v844f91;
assign v855002 = ENQ_p & v856553 | !ENQ_p & v85658a;
assign v857649 = ENQ_p & v86b41a | !ENQ_p & v8565c6;
assign v8541a9 = jx1_p & v856b69 | !jx1_p & v8a30d8;
assign v8a3354 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8567c7;
assign v855658 = jx2_p & v85ecbc | !jx2_p & v855386;
assign v855700 = RtoB_ACK1_p & v8556fc | !RtoB_ACK1_p & v876637;
assign v855acd = jx0_p & v8a3045 | !jx0_p & v8a2a91;
assign v8568b8 = ENQ_p & v856c57 | !ENQ_p & v8a3095;
assign v8552de = StoB_REQ0_p & v854b2f | !StoB_REQ0_p & v87d011;
assign v8a33af = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v856e7f;
assign v8a3339 = jx2_p & v856b4c | !jx2_p & v844f91;
assign v856467 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & !v8a2c94;
assign v8a2f1e = RtoB_ACK0_p & v8836e5 | !RtoB_ACK0_p & v856e02;
assign v855f89 = stateG7_1_p & v855ab2 | !stateG7_1_p & v855b5d;
assign v856639 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8a3036;
assign v856651 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8560c5;
assign v8a3233 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v854b1a;
assign v8559d2 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & v8553e7;
assign v8a30e5 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v867265;
assign v8a3156 = jx0_p & v8a32cc | !jx0_p & v855bae;
assign v8563c1 = jx0_p & v852505 | !jx0_p & v844f9d;
assign v854ff9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3265;
assign v844fad = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v8a314d = jx0_p & v85528e | !jx0_p & !v855ed8;
assign v855426 = jx0_p & v856aac | !jx0_p & v8562b9;
assign v8560e2 = ENQ_p & v8574ba | !ENQ_p & v855e7a;
assign v8a2faa = StoB_REQ1_p & v8549db | !StoB_REQ1_p & v8a31ff;
assign v855069 = RtoB_ACK0_p & v856e74 | !RtoB_ACK0_p & v856dec;
assign v857624 = jx1_p & v856982 | !jx1_p & v844f91;
assign v8a3395 = StoB_REQ1_p & v854bcd | !StoB_REQ1_p & v857452;
assign v854b5e = jx2_p & v8a31a2 | !jx2_p & v855254;
assign v870eb8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v8552c8 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v855eb2;
assign v855a8a = RtoB_ACK0_p & v854f1c | !RtoB_ACK0_p & v85682b;
assign v855d98 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a3269;
assign v855ac2 = EMPTY_p & v857aaa | !EMPTY_p & v8a2b13;
assign v856c11 = BtoR_REQ1_p & v857595 | !BtoR_REQ1_p & v8556a7;
assign v85768c = ENQ_p & v85741f | !ENQ_p & v855505;
assign v855505 = jx2_p & v844f91 | !jx2_p & v856b86;
assign v857775 = EMPTY_p & v8a30b5 | !EMPTY_p & v8a302d;
assign v86f7aa = EMPTY_p & v854f2f | !EMPTY_p & v8a30ec;
assign v8a30c7 = BtoS_ACK0_p & v85681c | !BtoS_ACK0_p & v8a326f;
assign v8a2b95 = jx0_p & v8578fc | !jx0_p & v855a8f;
assign v8a333f = ENQ_p & v8a324a | !ENQ_p & v856847;
assign v856432 = ENQ_p & v85413e | !ENQ_p & v844f91;
assign v8a29dc = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v8551dd;
assign v8a3287 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v888ec4;
assign v8a33d5 = BtoS_ACK0_p & v855311 | !BtoS_ACK0_p & v8a338c;
assign v8a30b6 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a3208;
assign v8a31b3 = BtoS_ACK0_p & v857880 | !BtoS_ACK0_p & !v8a3340;
assign v855850 = FULL_p & v85759c | !FULL_p & v8a30be;
assign v854ffe = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8558ad;
assign v8a2894 = ENQ_p & v8a302c | !ENQ_p & v844f91;
assign v8a2fd8 = ENQ_p & v86178d | !ENQ_p & v85660e;
assign v8569fe = ENQ_p & v8a324a | !ENQ_p & v8a2d44;
assign v86eb76 = jx1_p & v8a2dfa | !jx1_p & v85413e;
assign v8574ba = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v856705;
assign v8a2448 = jx0_p & v855858 | !jx0_p & !v855d6a;
assign v856443 = jx1_p & v85606a | !jx1_p & v8a3214;
assign v855418 = jx0_p & v8557e6 | !jx0_p & v856761;
assign v844f91 = 1;
assign v8a336b = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v855912;
assign v8a328d = BtoS_ACK0_p & v856883 | !BtoS_ACK0_p & v8550a0;
assign v8a336a = StoB_REQ0_p & v8a2b0e | !StoB_REQ0_p & v883709;
assign v88abb8 = jx0_p & v8a3289 | !jx0_p & !v8a3050;
assign v8a2f7a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8a2a8c;
assign v856543 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v854ee4;
assign v861d68 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86da55;
assign v8573b7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3112;
assign v8a3362 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8738b2;
assign v8a2f9b = BtoS_ACK0_p & v8a3379 | !BtoS_ACK0_p & v88ab71;
assign v8a31f6 = stateG12_p & v8574ba | !stateG12_p & v844f91;
assign v855709 = jx2_p & v8556c1 | !jx2_p & v8a31f2;
assign v8a3376 = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v873613;
assign v856723 = ENQ_p & v87c729 | !ENQ_p & v8a3160;
assign v856495 = stateG7_1_p & v856372 | !stateG7_1_p & v85ab38;
assign v8960ee = EMPTY_p & v8551da | !EMPTY_p & v8a330a;
assign v8a2d8d = BtoS_ACK0_p & v8564d2 | !BtoS_ACK0_p & v8557f6;
assign v877887 = StoB_REQ3_p & v8a312e | !StoB_REQ3_p & v844f91;
assign v855d3a = stateG7_1_p & v854c4e | !stateG7_1_p & v8a30c3;
assign v855564 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3184;
assign v85570e = jx2_p & v8a289a | !jx2_p & v85741f;
assign v855783 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f99;
assign v85759c = ENQ_p & v855f60 | !ENQ_p & v8a33c4;
assign v883759 = ENQ_p & v86b41a | !ENQ_p & v8a302f;
assign v854cad = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8561e7;
assign v85765d = jx1_p & v85ab66 | !jx1_p & v855268;
assign v854f9b = jx1_p & v854194 | !jx1_p & v85601a;
assign v85575f = jx0_p & v89fce5 | !jx0_p & v856b69;
assign v8a311c = StoB_REQ1_p & v8a3363 | !StoB_REQ1_p & v8a3101;
assign v85690e = jx2_p & v8558ea | !jx2_p & !v8578b4;
assign v868e49 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8532c4;
assign v854d3e = jx1_p & v85606a | !jx1_p & !v855418;
assign v85522d = StoB_REQ0_p & v85751a | !StoB_REQ0_p & v856075;
assign v86aa3d = EMPTY_p & v8553d5 | !EMPTY_p & v8a3182;
assign v867ef3 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v855ef6;
assign v856884 = EMPTY_p & v856b58 | !EMPTY_p & v8a3279;
assign BtoS_ACK3_n = !v86180e;
assign v855e00 = StoB_REQ4_p & v844fa0 | !StoB_REQ4_p & !v844f91;
assign v857543 = jx1_p & v856624 | !jx1_p & !v8a2448;
assign v8a30eb = BtoS_ACK0_p & v844fe7 | !BtoS_ACK0_p & v8a2b82;
assign v8579a9 = BtoS_ACK1_p & v8a3170 | !BtoS_ACK1_p & v856e34;
assign v856abb = jx1_p & v854b14 | !jx1_p & v844f91;
assign v85601a = jx0_p & v855011 | !jx0_p & v8550fb;
assign v8549ca = RtoB_ACK0_p & v8a3027 | !RtoB_ACK0_p & v8a31e3;
assign v856264 = BtoR_REQ1_p & v896174 | !BtoR_REQ1_p & v856bfd;
assign v8a3167 = jx2_p & v86f537 | !jx2_p & v857624;
assign v87532a = jx0_p & v8a3179 | !jx0_p & !v8a33de;
assign v8a33ac = jx1_p & v844f91 | !jx1_p & v8a3278;
assign v8a294c = BtoS_ACK2_p & v8a33c1 | !BtoS_ACK2_p & v8576bc;
assign v8a287f = stateG7_1_p & v8a322c | !stateG7_1_p & v856784;
assign v856e26 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8679b5;
assign v856041 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8a2dbf;
assign v856545 = jx1_p & v8a2fd5 | !jx1_p & v88abf3;
assign v85a4b3 = stateG12_p & v844f91 | !stateG12_p & !v8a3151;
assign v855531 = StoB_REQ1_p & v8630d3 | !StoB_REQ1_p & v89caa5;
assign v855600 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8630d3;
assign v8a3036 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v85523e;
assign v8a31ac = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v855d34;
assign v8a3077 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a33c2;
assign v855ba9 = jx1_p & v856624 | !jx1_p & !v855faf;
assign v8a31d5 = jx0_p & v86a9c5 | !jx0_p & v85606a;
assign v85581e = StoB_REQ3_p & v854c76 | !StoB_REQ3_p & v85523e;
assign v8a325b = StoB_REQ1_p & v8549db | !StoB_REQ1_p & v855d98;
assign v856b4c = jx1_p & v844f91 | !jx1_p & !v855221;
assign v8a3081 = BtoS_ACK4_p & v855e00 | !BtoS_ACK4_p & v844f9d;
assign v856c7e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3147;
assign v86c364 = StoB_REQ0_p & v855600 | !StoB_REQ0_p & v8a3116;
assign v8574ef = RtoB_ACK0_p & v854f98 | !RtoB_ACK0_p & v88abaa;
assign v856b86 = jx1_p & v855b6e | !jx1_p & v844f91;
assign v8563cf = ENQ_p & v857a8e | !ENQ_p & v8a32c3;
assign v85e22c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v87c759;
assign v855c86 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v85586d;
assign v8a2ef9 = RtoB_ACK1_p & v8554d7 | !RtoB_ACK1_p & v855218;
assign v855d5e = BtoS_ACK1_p & v856422 | !BtoS_ACK1_p & v857619;
assign v85a3c4 = EMPTY_p & v854a55 | !EMPTY_p & v8553df;
assign v8a2c28 = DEQ_p & v88ab6c | !DEQ_p & v8a329a;
assign v8a31cc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v856b2a;
assign v856313 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a3203;
assign v8a328b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85a3a7;
assign v8a3203 = StoB_REQ1_p & v8549db | !StoB_REQ1_p & v8a0e55;
assign v8a3197 = DEQ_p & v8551f9 | !DEQ_p & v8a331f;
assign v8a3270 = BtoS_ACK1_p & v8a333a | !BtoS_ACK1_p & v854fff;
assign v85544e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883cb2;
assign v8561a3 = jx2_p & v856195 | !jx2_p & v8579da;
assign v8a3275 = BtoS_ACK0_p & v855eb2 | !BtoS_ACK0_p & v85594d;
assign v8a313f = jx2_p & v854e8e | !jx2_p & !v855046;
assign v88ab9b = EMPTY_p & v8541c7 | !EMPTY_p & v8617c9;
assign v8a302e = jx2_p & v8a30a5 | !jx2_p & v844fa9;
assign v8a32f2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883cb1;
assign v8a2e42 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8a3220;
assign v856e0b = StoB_REQ1_p & v8a3130 | !StoB_REQ1_p & v856e10;
assign v855218 = EMPTY_p & v8a30af | !EMPTY_p & v8a2b13;
assign v855d84 = jx1_p & v8a2fd5 | !jx1_p & v85bce8;
assign v85be20 = jx0_p & v8a32c0 | !jx0_p & v8a2daf;
assign v86c421 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a33c1;
assign v8a2ef0 = ENQ_p & v85570e | !ENQ_p & v8a310e;
assign v8a317b = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v85509f;
assign v8a3329 = ENQ_p & v844f91 | !ENQ_p & v8a329f;
assign v888ec4 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a3080;
assign v8a3045 = BtoS_ACK0_p & v844fa0 | !BtoS_ACK0_p & v88ab87;
assign v856863 = BtoS_ACK1_p & v8a3032 | !BtoS_ACK1_p & v8a32ea;
assign v8565de = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v8555ef;
assign v8a30d8 = jx0_p & v8a30eb | !jx0_p & !v86aa28;
assign v85747f = jx0_p & v855a9b | !jx0_p & v844f91;
assign v8a3159 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8a2b16;
assign v8566d2 = jx0_p & v88ab9d | !jx0_p & !v8a24a6;
assign v8a3320 = BtoR_REQ1_p & v8a32e1 | !BtoR_REQ1_p & v8a32ef;
assign v85413e = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8573cd;
assign v856ac3 = jx1_p & v85606a | !jx1_p & !v8a31ba;
assign v8562e3 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v857b78;
assign v85adee = jx0_p & v8a2fa6 | !jx0_p & v854194;
assign v857866 = BtoS_ACK1_p & v854b7c | !BtoS_ACK1_p & !v8a3097;
assign v85756f = jx2_p & v855e0d | !jx2_p & v8579da;
assign v854ffa = stateG7_1_p & v8a3267 | !stateG7_1_p & v857674;
assign v8559e7 = jx2_p & v8a30e6 | !jx2_p & v85413e;
assign v8550b4 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86e4e3;
assign v8a3269 = StoB_REQ2_p & v856e2b | !StoB_REQ2_p & v8560ec;
assign v854f90 = StoB_REQ0_p & v8553e6 | !StoB_REQ0_p & v856b54;
assign v857b07 = StoB_REQ2_p & v85791e | !StoB_REQ2_p & v85be78;
assign v855bae = BtoS_ACK0_p & v857880 | !BtoS_ACK0_p & v8a338b;
assign v855735 = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v8a331c;
assign v8a32b6 = jx0_p & v8a330f | !jx0_p & !v8a3309;
assign v8711d9 = StoB_REQ3_p & v844f9d | !StoB_REQ3_p & v844f91;
assign v86aa4d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a33ce;
assign v876d41 = ENQ_p & v844fa9 | !ENQ_p & !v844f91;
assign v856c01 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a3389;
assign v85628f = jx0_p & v8a2a05 | !jx0_p & v8550fb;
assign v8541c7 = ENQ_p & v8574ba | !ENQ_p & v844f91;
assign v855d45 = jx0_p & v8a320f | !jx0_p & v8559aa;
assign v85ecbc = jx1_p & v8a3151 | !jx1_p & v85510d;
assign v8573a4 = jx0_p & v8a30b6 | !jx0_p & v85617a;
assign v88ab6c = ENQ_p & v8a324a | !ENQ_p & v85ecc8;
assign v88abd1 = DEQ_p & v855e0c | !DEQ_p & v856432;
assign v8a330c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855528;
assign v883cb8 = jx2_p & v8568ac | !jx2_p & v87c763;
assign v8a33c1 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v855b05;
assign v8a320e = stateG7_1_p & v8a30cd | !stateG7_1_p & v8a2bb4;
assign v854ae5 = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v856c23;
assign v854a89 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85ab2e;
assign v85ecc8 = jx2_p & v85a48b | !jx2_p & !v8a30e2;
assign v883756 = RtoB_ACK0_p & v856945 | !RtoB_ACK0_p & v8550af;
assign v8a2dfb = jx1_p & v8a2fba | !jx1_p & v8a329d;
assign v855674 = jx1_p & v888ed9 | !jx1_p & v85419c;
assign v896294 = EMPTY_p & v8a32bd | !EMPTY_p & !v854fc7;
assign v8a3128 = StoB_REQ2_p & v85532e | !StoB_REQ2_p & v872af1;
assign v85682b = stateG7_1_p & v8560a3 | !stateG7_1_p & v86179a;
assign v854d07 = DEQ_p & v8579f4 | !DEQ_p & v854a35;
assign v87e83a = jx2_p & v854d01 | !jx2_p & !v8a326b;
assign v8a3142 = jx2_p & v85778c | !jx2_p & !v8a317f;
assign v8552c6 = BtoS_ACK0_p & v85681c | !BtoS_ACK0_p & v8a330c;
assign v8a2d93 = BtoS_ACK2_p & v88b745 | !BtoS_ACK2_p & v8a3292;
assign v85646a = jx0_p & v8a3387 | !jx0_p & v856786;
assign v8a32e1 = RtoB_ACK0_p & v855db2 | !RtoB_ACK0_p & !v844f91;
assign v8555ef = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f99;
assign v869886 = StoB_REQ4_p & v8a2f21 | !StoB_REQ4_p & !v844f91;
assign v855c15 = RtoB_ACK1_p & v8a31e6 | !RtoB_ACK1_p & v8a3118;
assign v8a28d0 = EMPTY_p & v8a32c6 | !EMPTY_p & v8a3040;
assign BtoS_ACK0_n = v883775;
assign v8a303e = ENQ_p & v87c729 | !ENQ_p & v871174;
assign v88a46f = BtoR_REQ0_p & v8a3299 | !BtoR_REQ0_p & v8a3321;
assign v8961a6 = jx2_p & v86f537 | !jx2_p & v8a306b;
assign v8a32ba = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & !v856422;
assign BtoS_ACK5_n = !v86aa64;
assign v8a315d = StoB_REQ2_p & v8a308c | !StoB_REQ2_p & !v844f91;
assign v8836e5 = EMPTY_p & v8a2837 | !EMPTY_p & v854d1f;
assign v8961a7 = DEQ_p & v8551f9 | !DEQ_p & v856b8f;
assign v856b13 = stateG7_1_p & v855c15 | !stateG7_1_p & v8a3118;
assign v8a30de = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v855f43;
assign v856352 = BtoS_ACK2_p & v8567ec | !BtoS_ACK2_p & v8a2485;
assign v85a071 = jx0_p & v8a30e7 | !jx0_p & !v8a2fd5;
assign v856553 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fab;
assign v8557a6 = BtoS_ACK0_p & v8a30f6 | !BtoS_ACK0_p & v8a3272;
assign v8a3304 = DEQ_p & v8563cf | !DEQ_p & v8a2f08;
assign v8a339b = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8a3269;
assign v85635c = StoB_REQ4_p & v8a336c | !StoB_REQ4_p & !v844f91;
assign v8a3225 = BtoS_ACK1_p & v854a11 | !BtoS_ACK1_p & v8566ad;
assign v8a2cc7 = ENQ_p & v856553 | !ENQ_p & !v855b2c;
assign v8a3333 = ENQ_p & v8574ba | !ENQ_p & v854eff;
assign v854fcb = ENQ_p & v85610f | !ENQ_p & v8a33a5;
assign v856982 = jx0_p & v857b70 | !jx0_p & v844f91;
assign v88ea49 = BtoR_REQ0_p & v8a28a9 | !BtoR_REQ0_p & !v8a3320;
assign v854f52 = BtoS_ACK4_p & v8573ee | !BtoS_ACK4_p & v8a2f21;
assign v8a32e8 = ENQ_p & v844f91 | !ENQ_p & v8a3339;
assign v8a3356 = BtoS_ACK2_p & v8711d9 | !BtoS_ACK2_p & v856e7f;
assign v8a333a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v88b745;
assign v855b1d = EMPTY_p & v883759 | !EMPTY_p & v8a302d;
assign v85659e = jx1_p & v844f91 | !jx1_p & v8541e6;
assign v8a3099 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3144;
assign v8558e6 = BtoS_ACK0_p & v8a30f6 | !BtoS_ACK0_p & v856799;
assign v8561e7 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854a17;
assign v8a3228 = RtoB_ACK1_p & v8559bc | !RtoB_ACK1_p & v855ea7;
assign v8a3336 = BtoS_ACK1_p & v8a333a | !BtoS_ACK1_p & v8a31b6;
assign v8a2c17 = jx1_p & v85606a | !jx1_p & !v8a30ba;
assign v8a30f7 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a3175;
assign v8551da = ENQ_p & v8a324a | !ENQ_p & v8549fe;
assign v8a30b4 = StoB_REQ0_p & v8a30b3 | !StoB_REQ0_p & v857866;
assign v8a3154 = jx2_p & v8a29cd | !jx2_p & !v855df9;
assign v856176 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v855783;
assign v8558ad = BtoS_ACK1_p & v854a11 | !BtoS_ACK1_p & v8a3140;
assign v86c9ca = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a294c;
assign v8a283f = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a24df;
assign v8573cd = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a3314;
assign v8a2c94 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8a3350;
assign v8a3367 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v855bf8;
assign v867265 = StoB_REQ1_p & v854c82 | !StoB_REQ1_p & v8a2ae0;
assign v854138 = jx0_p & v8a3260 | !jx0_p & !v857a21;
assign v856d89 = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & v8685f8;
assign v8a3131 = EMPTY_p & v8a329c | !EMPTY_p & v854a07;
assign v858911 = jx1_p & v844f91 | !jx1_p & v85a4b2;
assign v85525c = jx2_p & v854cd0 | !jx2_p & !v8a304d;
assign v86aa63 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f9d;
assign v8a31bc = DEQ_p & v883741 | !DEQ_p & v854994;
assign v857619 = StoB_REQ1_p & v8555ef | !StoB_REQ1_p & v857785;
assign v8a3293 = EMPTY_p & v8541c7 | !EMPTY_p & v85a4b4;
assign v8a2ec1 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v855eb3;
assign v857694 = jx2_p & v89612f | !jx2_p & !v8a30bf;
assign v8a2972 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v844f91;
assign v8a2bfa = jx2_p & v8a3261 | !jx2_p & !v85685d;
assign v8a3083 = ENQ_p & v855f60 | !ENQ_p & v8a32ae;
assign v8a30e6 = jx1_p & v855565 | !jx1_p & v85413e;
assign v8a31d1 = jx0_p & v8a2fb0 | !jx0_p & v8a2d8d;
assign v8a291b = EMPTY_p & v8a2837 | !EMPTY_p & v8a3066;
assign v854d20 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a31bd;
assign v8551f9 = ENQ_p & v855653 | !ENQ_p & v86fe32;
assign v855ef6 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9b;
assign v8a319c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a33b3;
assign v8558fa = ENQ_p & v85741f | !ENQ_p & v8a30ef;
assign v8a32d3 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a2b63;
assign v8568ac = jx1_p & v856b69 | !jx1_p & v857a4d;
assign v883cae = RtoB_ACK1_p & v8a291b | !RtoB_ACK1_p & v861800;
assign v873853 = RtoB_ACK1_p & v8a0e4e | !RtoB_ACK1_p & v854fe3;
assign v8a321e = jx2_p & v8a29d0 | !jx2_p & !v85685d;
assign v855011 = BtoS_ACK0_p & v87c725 | !BtoS_ACK0_p & v85522b;
assign v855ae0 = ENQ_p & v8575b5 | !ENQ_p & v8a2e43;
assign v896106 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v877670;
assign v855957 = RtoB_ACK0_p & v8a3187 | !RtoB_ACK0_p & v85554e;
assign v8a2fba = BtoS_ACK0_p & v8a3089 | !BtoS_ACK0_p & v85e22c;
assign v8691ce = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3054;
assign v856d52 = jx1_p & v85499f | !jx1_p & !v856023;
assign v85a3a3 = EMPTY_p & v856432 | !EMPTY_p & v85562c;
assign v8a3179 = BtoS_ACK0_p & v8a2972 | !BtoS_ACK0_p & v8a3075;
assign v8a33da = BtoS_ACK0_p & v854b7c | !BtoS_ACK0_p & v8a30b4;
assign v8558ec = BtoS_ACK0_p & v8a2972 | !BtoS_ACK0_p & v854b6c;
assign v8a24df = BtoS_ACK4_p & v854ee4 | !BtoS_ACK4_p & v8685f8;
assign v8a3360 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85621e;
assign v866b88 = ENQ_p & v8a32da | !ENQ_p & !v844f91;
assign v8567b5 = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v855078;
assign v8a326c = ENQ_p & v8a3142 | !ENQ_p & v8a329f;
assign v8a29f8 = jx1_p & v855d7a | !jx1_p & !v855b2d;
assign v856a98 = jx2_p & v857aee | !jx2_p & v8a3090;
assign v855bc8 = jx0_p & v856aac | !jx0_p & !v8562b9;
assign v8a2d1f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855735;
assign v8a2e9b = StoB_REQ2_p & v856acb | !StoB_REQ2_p & v8a3217;
assign v8a3241 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v88b745;
assign v855791 = StoB_REQ0_p & v8a2893 | !StoB_REQ0_p & v8a313d;
assign v855edf = StoB_REQ0_p & v8550f3 | !StoB_REQ0_p & v844f91;
assign v854eb2 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a33ec;
assign v8a3214 = jx0_p & v85663b | !jx0_p & v855879;
assign v854a0a = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a302a;
assign v8a2c75 = jx2_p & v854c99 | !jx2_p & !v85793b;
assign v855042 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v855833;
assign v873869 = StoB_REQ1_p & v8555ef | !StoB_REQ1_p & !v8551d0;
assign v8a28b9 = StoB_REQ2_p & v883730 | !StoB_REQ2_p & v8960f3;
assign v8a30fe = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v854e55;
assign v8561e1 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v855eb2;
assign v8574f8 = jx2_p & v8a33ac | !jx2_p & !v8a2cbd;
assign v857674 = EMPTY_p & v8560e2 | !EMPTY_p & v8962fa;
assign v8554f7 = stateG12_p & v856553 | !stateG12_p & v844f91;
assign v8a3318 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v89625f;
assign v856903 = jx0_p & v856653 | !jx0_p & !v844f91;
assign v8a315a = jx0_p & v8a3046 | !jx0_p & v854194;
assign v8a31fa = jx1_p & v844f91 | !jx1_p & !v88abb8;
assign v85607f = jx0_p & v8550e8 | !jx0_p & v8a3275;
assign v8a318e = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8a283f;
assign v85675f = StoB_REQ1_p & v8a3356 | !StoB_REQ1_p & v8a33af;
assign v855533 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a2e94;
assign v8a320a = jx0_p & v8562f8 | !jx0_p & v8a2d8d;
assign v8560bc = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v8551d0;
assign v8549e6 = jx2_p & v8a2d10 | !jx2_p & v8a2d94;
assign v854f04 = jx2_p & v8a3300 | !jx2_p & v8565a7;
assign v855786 = ENQ_p & v85741f | !ENQ_p & v8561a3;
assign v856349 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a339d;
assign v8558ea = jx1_p & v85606a | !jx1_p & v855631;
assign v87c6f7 = RtoB_ACK1_p & v854988 | !RtoB_ACK1_p & v85531c;
assign v8a2d29 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8a2c6c;
assign v857a0d = stateG7_1_p & v8a33be | !stateG7_1_p & v844f91;
assign v8a31a9 = EMPTY_p & v857487 | !EMPTY_p & v8a3197;
assign v8a3261 = jx1_p & v854194 | !jx1_p & v8a2b95;
assign v8a30c9 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8555ef;
assign v888ecd = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a2c6b;
assign v855912 = StoB_REQ0_p & v86a9cb | !StoB_REQ0_p & v8567b8;
assign v8a3149 = RtoB_ACK1_p & v856884 | !RtoB_ACK1_p & v855414;
assign v8a307d = jx1_p & v844f91 | !jx1_p & v85628f;
assign v855583 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8555d3;
assign v854e78 = StoB_REQ0_p & v8a30f7 | !StoB_REQ0_p & v844f91;
assign v8a3022 = EMPTY_p & v855c80 | !EMPTY_p & v855283;
assign v85aaf7 = jx1_p & v8a2fba | !jx1_p & v8a2a54;
assign v85746e = jx1_p & v844f91 | !jx1_p & !v8a31b0;
assign v8960f3 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v85635c;
assign v854a11 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9d;
assign v8a3030 = jx2_p & v8654fb | !jx2_p & !v8a30e2;
assign v8a0e3c = jx1_p & v844f91 | !jx1_p & !v871154;
assign v8567ec = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v85523e;
assign v8a3185 = DEQ_p & v8a3038 | !DEQ_p & v8a313e;
assign v855941 = jx0_p & v8560fa | !jx0_p & v8a3376;
assign v870ea9 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v854d20;
assign v85743a = ENQ_p & v8a2a7f | !ENQ_p & !v8a33c0;
assign v8557f8 = RtoB_ACK0_p & v854c39 | !RtoB_ACK0_p & v8a33e5;
assign v8a2e94 = StoB_REQ1_p & v88a44b | !StoB_REQ1_p & v844f91;
assign v8a33aa = jx1_p & v844f91 | !jx1_p & v8557e1;
assign v85745e = jx1_p & v85a4b3 | !jx1_p & v844f91;
assign v88abf3 = jx0_p & v8738de | !jx0_p & v8a3273;
assign v856ad2 = stateG7_1_p & v85555f | !stateG7_1_p & v8573a2;
assign v88abc5 = EMPTY_p & v8554b2 | !EMPTY_p & v855fb5;
assign v85678b = DEQ_p & v855f95 | !DEQ_p & v8a330a;
assign v855bf8 = RtoB_ACK0_p & v857a0d | !RtoB_ACK0_p & v8a2fa9;
assign v8a3170 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8567ec;
assign v8a327a = jx0_p & v855858 | !jx0_p & !v854b8e;
assign v8a33e5 = stateG7_1_p & v8a3346 | !stateG7_1_p & v8a2b29;
assign v855e7a = jx2_p & v8549bd | !jx2_p & !v8a3200;
assign v871675 = BtoS_ACK1_p & v844fa0 | !BtoS_ACK1_p & v856af3;
assign v8a2ce0 = jx1_p & v856786 | !jx1_p & v8551a3;
assign v8a31b5 = stateG7_1_p & v8a3173 | !stateG7_1_p & v8a31df;
assign v857418 = jx2_p & v8a2ce0 | !jx2_p & !v85793b;
assign v85540d = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9b;
assign v8a3183 = jx0_p & v85528e | !jx0_p & !v871138;
assign v8a30bf = jx1_p & v8a3158 | !jx1_p & v856cee;
assign v854d1f = DEQ_p & v8a2ef0 | !DEQ_p & v856535;
assign v8a2e77 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a287d;
assign v856288 = jx0_p & v8a29ad | !jx0_p & !v8a3235;
assign v8a3193 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v85586d;
assign v8a2b0e = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8a3377;
assign v855221 = jx0_p & v8a30e9 | !jx0_p & !v844f91;
assign v855ce1 = stateG7_1_p & v8a31a9 | !stateG7_1_p & v8a309e;
assign v85e7e0 = jx1_p & v844f91 | !jx1_p & v8617f7;
assign v8a3260 = BtoS_ACK0_p & v857a31 | !BtoS_ACK0_p & v855748;
assign v854e55 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8a315d;
assign v854c40 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & v854a71;
assign v854edc = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8559ce;
assign v8a31cd = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v855583;
assign v88372d = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v855ef6;
assign v8a30c2 = StoB_REQ3_p & v8685f8 | !StoB_REQ3_p & v844f91;
assign v856575 = jx1_p & v844f91 | !jx1_p & !v856df4;
assign v8a3046 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8550b4;
assign v8573a2 = EMPTY_p & v8a3155 | !EMPTY_p & !v8a2891;
assign v8a31ea = jx1_p & v8a32b6 | !jx1_p & v85509e;
assign v855d70 = DEQ_p & v8a3286 | !DEQ_p & v8a296b;
assign v854f97 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v855ee6;
assign v86da55 = BtoS_ACK1_p & v8a2972 | !BtoS_ACK1_p & v856c7e;
assign v854988 = EMPTY_p & v8a3202 | !EMPTY_p & !v8a2891;
assign v8a309a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a3033;
assign v861796 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844faf;
assign v8a30a3 = jx2_p & v8a33aa | !jx2_p & v844f91;
assign v8a32bd = ENQ_p & v85610f | !ENQ_p & v8a3167;
assign v85eb9f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v855783;
assign v854fc1 = ENQ_p & v8549e6 | !ENQ_p & v86cbc9;
assign v8738b2 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v856ad7;
assign v8a337f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856422;
assign v8550f3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v856111;
assign v8a0dfa = jx1_p & v85be20 | !jx1_p & v854cc4;
assign v8a3272 = StoB_REQ0_p & v85eb80 | !StoB_REQ0_p & v85634e;
assign v856441 = BtoS_ACK0_p & v855eb2 | !BtoS_ACK0_p & v8562af;
assign v855137 = DEQ_p & v85798c | !DEQ_p & v8a2ff2;
assign v856847 = jx2_p & v8560ff | !jx2_p & !v8a31ea;
assign v8962ff = BtoR_REQ0_p & v844fa1 | !BtoR_REQ0_p & v8a3367;
assign v85aad7 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v857b07;
assign v8a32a9 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v8a3193;
assign v8a31aa = jx0_p & v8a2fb0 | !jx0_p & v844f91;
assign v856730 = ENQ_p & v85610f | !ENQ_p & v8961a6;
assign v8a3075 = StoB_REQ0_p & v854b2f | !StoB_REQ0_p & v8a321c;
assign v856d91 = ENQ_p & v844fa9 | !ENQ_p & !v854aa0;
assign v854fe3 = EMPTY_p & v85d977 | !EMPTY_p & v8961a7;
assign v855ebf = EMPTY_p & v8a3079 | !EMPTY_p & v8567aa;
assign v8a327f = jx2_p & v8a307d | !jx2_p & !v8a3200;
assign v8a3372 = jx0_p & v855858 | !jx0_p & !v856624;
assign v855e27 = stateG7_1_p & v8a24c7 | !stateG7_1_p & v883754;
assign v8a336e = FULL_p & v8a331f | !FULL_p & v85683b;
assign v854c4e = EMPTY_p & v8a303e | !EMPTY_p & v854cf3;
assign v8579cf = jx1_p & v8a3151 | !jx1_p & v854138;
assign v8567b8 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v855c5f;
assign v8578fc = BtoS_ACK0_p & v87c725 | !BtoS_ACK0_p & v8a32f2;
assign v8a31b0 = jx0_p & v855894 | !jx0_p & !v8566e1;
assign v8565ba = jx2_p & v855681 | !jx2_p & v85765d;
assign v854b33 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v854bcd;
assign v8662d9 = EMPTY_p & v8a282b | !EMPTY_p & v8567aa;
assign DEQ_n = !v88ea49;
assign v856e5f = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8a2e4a;
assign v856302 = StoB_REQ3_p & v8560ea | !StoB_REQ3_p & v844fb1;
assign v8a3392 = jx0_p & v8579f3 | !jx0_p & v8a3361;
assign v8559aa = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v855df1;
assign v8a3415 = jx0_p & v89626e | !jx0_p & v844f91;
assign v8a3070 = jx1_p & v844f91 | !jx1_p & v8a2479;
assign v856b54 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8551c8;
assign v8a33ec = StoB_REQ1_p & v8549db | !StoB_REQ1_p & v8a339b;
assign v8a3200 = jx1_p & v8a33ad | !jx1_p & !v854194;
assign v8550db = RtoB_ACK0_p & v856ad2 | !RtoB_ACK0_p & v8a31b5;
assign v856c9f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85540d;
assign v855748 = StoB_REQ0_p & v854b2f | !StoB_REQ0_p & v8a31b7;
assign v87c725 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a3086;
assign v85ec27 = jx1_p & v856b69 | !jx1_p & v8a335b;
assign v8a2a05 = BtoS_ACK0_p & v87c725 | !BtoS_ACK0_p & v85416e;
assign v857a91 = jx1_p & v8a33e8 | !jx1_p & v8574ba;
assign v8a284d = jx0_p & v8a30b3 | !jx0_p & v8a2fd5;
assign v855c79 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v8711c0;
assign v86aa4b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v856d89;
assign v8a30b8 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a3334;
assign v87bbfb = jx2_p & v873280 | !jx2_p & !v8a2eb6;
assign v844fe7 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a3170;
assign v8a3388 = jx0_p & v844f91 | !jx0_p & v8a2fd5;
assign v8a31af = ENQ_p & v8574eb | !ENQ_p & v8a304c;
assign v856c57 = jx2_p & v8567a3 | !jx2_p & !v8a326b;
assign v8a3284 = jx0_p & v8a3196 | !jx0_p & v88a469;
assign v8a307b = ENQ_p & v85413e | !ENQ_p & v8a30aa;
assign v8a29cd = jx1_p & v844f91 | !jx1_p & !v8a300d;
assign v855ead = ENQ_p & v8574ba | !ENQ_p & v8a2bfa;
assign v8a2a74 = BtoS_ACK0_p & v8a3129 | !BtoS_ACK0_p & v8a328a;
assign v8a323e = jx1_p & v85606a | !jx1_p & !v8a3242;
assign v856417 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a2ffa;
assign v8556fc = EMPTY_p & v85548d | !EMPTY_p & v857689;
assign v8961ac = jx0_p & v8962e0 | !jx0_p & v8a30c9;
assign v8a3108 = jx1_p & v8a2fba | !jx1_p & v85607f;
assign v8a305b = jx2_p & v8579cf | !jx2_p & v855df9;
assign v8553d5 = ENQ_p & v844f91 | !ENQ_p & !v8575a5;
assign v855e0e = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v869f3f;
assign v8575aa = ENQ_p & v8a3342 | !ENQ_p & v844f91;
assign v855935 = jx2_p & v854f9b | !jx2_p & !v855edc;
assign v8552f8 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v854188;
assign v8a329b = jx1_p & v844f91 | !jx1_p & !v8a2d5b;
assign v8a3223 = RtoB_ACK0_p & v8a33b1 | !RtoB_ACK0_p & v857a65;
assign v86a9e8 = EMPTY_p & v8568be | !EMPTY_p & v855d70;
assign v8550be = jx0_p & v85edf0 | !jx0_p & v855879;
assign v85eae9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8562e3;
assign v8a32a3 = BtoS_ACK0_p & v8561e1 | !BtoS_ACK0_p & v8a3253;
assign v86624f = jx0_p & v8a33da | !jx0_p & !v8a3151;
assign v855d54 = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v8a325b;
assign v8a329a = ENQ_p & v8a313f | !ENQ_p & v85ecc8;
assign v85791e = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v854f52;
assign v85500c = RtoB_ACK1_p & v88abc3 | !RtoB_ACK1_p & v8a3131;
assign v856737 = BtoR_REQ1_p & v85648f | !BtoR_REQ1_p & !v883756;
assign v8558d6 = jx0_p & v855894 | !jx0_p & v844f91;
assign v855b6e = jx0_p & v844f91 | !jx0_p & !v871138;
assign v8a3358 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v856731;
assign v855361 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v855311;
assign v856197 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a2e77;
assign v857b78 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a3350;
assign v8a33c7 = StoB_REQ1_p & v86f89c | !StoB_REQ1_p & v8a2e89;
assign v896289 = ENQ_p & v8a332a | !ENQ_p & !v8a338f;
assign v8a0e03 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v85523e;
assign v855b24 = ENQ_p & v8a324a | !ENQ_p & v854a8f;
assign v87c763 = jx1_p & v8a3031 | !jx1_p & v8a3181;
assign v854ccd = FULL_p & v854a55 | !FULL_p & v85768c;
assign v844fa9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v859301 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8a30b4;
assign v85677d = StoB_REQ0_p & v8a2f07 | !StoB_REQ0_p & v855cd9;
assign v8a3313 = jx0_p & v8a3098 | !jx0_p & v8a0de9;
assign v85576e = BtoS_ACK1_p & v854a11 | !BtoS_ACK1_p & v87116b;
assign v8a305e = BtoR_REQ1_p & v8a2f1e | !BtoR_REQ1_p & v855fec;
assign v854f8b = jx0_p & v8a2a74 | !jx0_p & v8a0de9;
assign v8654fb = jx1_p & v844f91 | !jx1_p & !v8a3153;
assign v857af8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a337e;
assign v85778e = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8558fe;
assign v857727 = EMPTY_p & v8a3243 | !EMPTY_p & !v8a31bc;
assign v857a65 = stateG7_1_p & v855e5a | !stateG7_1_p & v85a3a3;
assign v855ff1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854f20;
assign v85601f = ENQ_p & v8574eb | !ENQ_p & v857694;
assign v8553df = DEQ_p & v8575aa | !DEQ_p & v854a55;
assign v855eb3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855c6b;
assign v8a33cf = StoB_REQ0_p & v85614f | !StoB_REQ0_p & v855185;
assign v855858 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v854b2f;
assign v8a2f17 = ENQ_p & v8a324a | !ENQ_p & v8a32b8;
assign v8a33e8 = stateG12_p & v8574ba | !stateG12_p & v854194;
assign v8a30e1 = DEQ_p & v8575aa | !DEQ_p & v85768c;
assign v8a33a5 = jx2_p & v86f537 | !jx2_p & v856abb;
assign v883775 = BtoR_REQ0_p & v8a312d | !BtoR_REQ0_p & v856db6;
assign v8a3175 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8a29a5;
assign v8a33bc = RtoB_ACK1_p & v855845 | !RtoB_ACK1_p & v85a3c4;
assign v856799 = StoB_REQ0_p & v85778e | !StoB_REQ0_p & v8a3322;
assign v854a53 = BtoS_ACK1_p & v8a333a | !BtoS_ACK1_p & v87116a;
assign v856026 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8541c6;
assign jx2_n = !v888edb;
assign v85565b = stateG12_p & v855254 | !stateG12_p & v856624;
assign v8a306f = BtoS_ACK1_p & v88b745 | !BtoS_ACK1_p & v857534;
assign v856731 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a2e00;
assign v855cd9 = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v8a311c;
assign v856761 = BtoS_ACK0_p & v8711cf | !BtoS_ACK0_p & v856102;
assign v86d760 = RtoB_ACK0_p & v8a3293 | !RtoB_ACK0_p & v8a31cb;
assign v860488 = jx1_p & v85698e | !jx1_p & !v8579c7;
assign v88a458 = StoB_REQ1_p & v867273 | !StoB_REQ1_p & v855564;
assign v8a310e = jx2_p & v86917e | !jx2_p & v8579da;
assign v8566bd = jx2_p & v844f91 | !jx2_p & !v8a3381;
assign v8554b2 = ENQ_p & v856553 | !ENQ_p & !v86007c;
assign v8a31e5 = DEQ_p & v85a137 | !DEQ_p & v8a329a;
assign v8a306e = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v85ab2a;
assign v8574eb = jx2_p & v856ac3 | !jx2_p & v85765d;
assign v854e7c = StoB_REQ2_p & v856543 | !StoB_REQ2_p & v844f91;
assign v85640f = ENQ_p & v844f91 | !ENQ_p & v8a30d1;
assign v86e4e3 = BtoS_ACK1_p & v8a3186 | !BtoS_ACK1_p & v8a31fe;
assign v856be3 = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v88b745;
assign v855014 = BtoS_ACK0_p & v844fe7 | !BtoS_ACK0_p & v856e7b;
assign v8a31a2 = jx1_p & v8a3106 | !jx1_p & v855254;
assign v8573d3 = jx0_p & v859301 | !jx0_p & v8a3151;
assign v854d33 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & !v855c3e;
assign v855c9e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v856262;
assign v85ab66 = jx0_p & v8a32a7 | !jx0_p & v8557b8;
assign v854a8f = jx2_p & v863beb | !jx2_p & !v8a31ea;
assign v855d3e = RtoB_ACK0_p & v88abc5 | !RtoB_ACK0_p & v855f89;
assign v873fa6 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85509b;
assign v85ab14 = DEQ_p & v855fb0 | !DEQ_p & v8a3294;
assign v8a2be7 = stateG7_1_p & v854aed | !stateG7_1_p & v844f91;
assign v855db1 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v86aa63;
assign v856111 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & !v855ef6;
assign v8a32b9 = BtoS_ACK0_p & v8a3379 | !BtoS_ACK0_p & v856436;
assign v8a315e = jx0_p & v8a32df | !jx0_p & v85676f;
assign v8a0e17 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856543;
assign v856d80 = EMPTY_p & v88ab43 | !EMPTY_p & v8a3185;
assign v857a8e = jx2_p & v857a91 | !jx2_p & v8574ba;
assign v855e79 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87d033;
assign v8a3397 = EMPTY_p & v8a3333 | !EMPTY_p & v8962fa;
assign v8a31f2 = jx1_p & v855941 | !jx1_p & v856e47;
assign v8a3243 = ENQ_p & v856c57 | !ENQ_p & v88371a;
assign v854a35 = FULL_p & v856535 | !FULL_p & v855786;
assign v85ed6f = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v8711d9;
assign v8a30a6 = ENQ_p & v8559e7 | !ENQ_p & v844f91;
assign v8a3152 = BtoS_ACK0_p & v855311 | !BtoS_ACK0_p & !v856651;
assign v8a321d = BtoS_ACK0_p & v85ed6f | !BtoS_ACK0_p & v854ae3;
assign v856535 = ENQ_p & v85741f | !ENQ_p & v85756f;
assign v8a32cb = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8a30c2;
assign v854194 = BtoS_ACK0_p & v85681c | !BtoS_ACK0_p & v8550b4;
assign v8560aa = StoB_REQ0_p & v8a2f46 | !StoB_REQ0_p & v8a30bd;
assign v844fa0 = StoB_REQ5_n & v844f91 | !StoB_REQ5_n & !v844f91;
assign v85606a = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v8a338c;
assign v865fb9 = BtoS_ACK2_p & v8a3036 | !BtoS_ACK2_p & v8a2a3d;
assign v855681 = jx1_p & v85524b | !jx1_p & !v8a31ba;
assign v88375a = jx2_p & v8a3317 | !jx2_p & v8a2d94;
assign v86aa28 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8a2b0e;
assign v8a3334 = StoB_REQ2_p & v855ef6 | !StoB_REQ2_p & v8a32ba;
assign v8a32fd = StoB_REQ0_p & v85778e | !StoB_REQ0_p & v856467;
assign v8a3302 = RtoB_ACK1_p & v8a3187 | !RtoB_ACK1_p & v8711bb;
assign v855b2d = jx0_p & v855d2c | !jx0_p & !v8a2fba;
assign v8a2dc2 = StoB_REQ0_p & v8565de | !StoB_REQ0_p & v8a3330;
assign v8a24c7 = EMPTY_p & v855e06 | !EMPTY_p & v8a31e5;
assign v8a3379 = StoB_REQ1_p & v844f9f | !StoB_REQ1_p & v856639;
assign v8a319e = EMPTY_p & v85aab4 | !EMPTY_p & v8a327e;
assign v856678 = StoB_REQ0_p & v8a2b0e | !StoB_REQ0_p & v844f91;
assign v8a30c3 = EMPTY_p & v8a3221 | !EMPTY_p & v854cf3;
assign v8961ce = jx0_p & v8a0e4f | !jx0_p & v870eb8;
assign v855a47 = EMPTY_p & v855c80 | !EMPTY_p & v854204;
assign v855268 = jx0_p & v8a33d5 | !jx0_p & v85606a;
assign v8558ef = RtoB_ACK0_p & v8a288c | !RtoB_ACK0_p & v8a32d8;
assign v8a2a54 = jx0_p & v8558ec | !jx0_p & v8a3327;
assign v8a2ffa = BtoS_ACK1_p & v8a2972 | !BtoS_ACK1_p & v8a2bf7;
assign v888ed9 = jx0_p & v856c72 | !jx0_p & !v8a31fb;
assign v8961a8 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a322d;
assign v85531b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v857866;
assign v855a8f = BtoS_ACK0_p & v8a3246 | !BtoS_ACK0_p & v8691ce;
assign v85528a = jx2_p & v844f91 | !jx2_p & v85665d;
assign v85665d = jx1_p & v844f91 | !jx1_p & v8a3388;
assign v856256 = RtoB_ACK0_p & v855d3a | !RtoB_ACK0_p & v8a309d;
assign v8a30f0 = jx2_p & v855c77 | !jx2_p & v856b69;
assign v8a331a = RtoB_ACK1_p & v854b24 | !RtoB_ACK1_p & v86a9e8;
assign v8a2ff0 = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v8a33df;
assign v85660e = jx2_p & v856443 | !jx2_p & !v8a30ce;
assign v876d51 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9f;
assign v855a61 = DEQ_p & v866b88 | !DEQ_p & v8a2c6e;
assign v876637 = EMPTY_p & v85548d | !EMPTY_p & v8563d8;
assign v8a3096 = BtoS_ACK2_p & v8711d9 | !BtoS_ACK2_p & !v854ed3;
assign v844fc1 = stateG12_p & v844f91 | !stateG12_p & !v844f91;
assign v8a31fd = RtoB_ACK0_p & v856495 | !RtoB_ACK0_p & v86e908;
assign v8a3325 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8554bf;
assign v8557e6 = BtoS_ACK0_p & v855c79 | !BtoS_ACK0_p & v855791;
assign v87734d = FULL_p & v844f91 | !FULL_p & v8a2d0e;
assign v8a31b7 = BtoS_ACK1_p & v854b1e | !BtoS_ACK1_p & v857421;
assign v8a33b1 = EMPTY_p & v856432 | !EMPTY_p & v855fac;
assign v857595 = EMPTY_p & v856730 | !EMPTY_p & !v854fc7;
assign v844fab = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v857880 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v855311;
assign v8a32a6 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v857469;
assign v8a3132 = BtoS_ACK2_p & v844fa0 | !BtoS_ACK2_p & v85eda6;
assign v855185 = BtoS_ACK1_p & v8a3170 | !BtoS_ACK1_p & v85644e;
assign v8a326b = jx1_p & v8a3043 | !jx1_p & v8a3150;
assign v8567a3 = jx1_p & v844f91 | !jx1_p & v8a2fac;
assign v855c38 = EMPTY_p & v85601f | !EMPTY_p & v857689;
assign v8a31d8 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v855783;
assign v8a3032 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v856422;
assign v8563d8 = DEQ_p & v8a338e | !DEQ_p & v855850;
assign v8a32c3 = jx2_p & v85520c | !jx2_p & !v8a3200;
assign v8a31ba = jx0_p & v854feb | !jx0_p & v88abed;
assign v85ed1a = jx1_p & v856786 | !jx1_p & v8a3214;
assign v8a3062 = DEQ_p & v85743a | !DEQ_p & v85504a;
assign v8a0e69 = BtoR_REQ0_p & v855a8a | !BtoR_REQ0_p & v8a305e;
assign v8a30b3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v87c747 = stateG7_1_p & v8a3149 | !stateG7_1_p & v854fe3;
assign v855a6a = DEQ_p & v8563cf | !DEQ_p & v8a339f;
assign v855c3e = StoB_REQ3_p & v85635c | !StoB_REQ3_p & !v85523e;
assign v8a3286 = ENQ_p & v8a2a7f | !ENQ_p & !v8a305b;
assign v8a3202 = ENQ_p & v87e83a | !ENQ_p & v8a3095;
assign v8550c7 = EMPTY_p & v8564e9 | !EMPTY_p & v8a327e;
assign v8555d3 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8a24df;
assign v8a3198 = DEQ_p & v8a30a6 | !DEQ_p & v8a307b;
assign v856653 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8550f3;
assign v8a3048 = ENQ_p & v8574ba | !ENQ_p & v8566bd;
assign v85edf1 = BtoR_REQ0_p & v855d3e | !BtoR_REQ0_p & v85554c;
assign v8a2aed = StoB_REQ2_p & v8a33d3 | !StoB_REQ2_p & v8a32cb;
assign v8a30f8 = RtoB_ACK1_p & v855db2 | !RtoB_ACK1_p & !v844f91;
assign v8a306b = jx1_p & v883733 | !jx1_p & v844f91;
assign v856784 = EMPTY_p & v8a310d | !EMPTY_p & v855182;
assign v871138 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8565de;
assign v85a48b = jx1_p & v844f91 | !jx1_p & !v8566d2;
assign v8564d2 = StoB_REQ1_p & v8a333a | !StoB_REQ1_p & v844f91;
assign v8a320d = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v86f804;
assign v8a2a7f = jx2_p & v85745e | !jx2_p & v844f91;
assign v854994 = ENQ_p & v856aa1 | !ENQ_p & v856489;
assign v85ed68 = jx0_p & v856653 | !jx0_p & v871138;
assign v8a339a = StoB_REQ1_p & v873fa6 | !StoB_REQ1_p & v870eba;
assign v86178d = jx2_p & v8a2c17 | !jx2_p & v85765d;
assign v8a3207 = StoB_REQ0_p & v85778e | !StoB_REQ0_p & v844f91;
assign v8a29a5 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v856d89;
assign v8a329d = jx0_p & v89626e | !jx0_p & v856441;
assign v8549bd = jx1_p & v854194 | !jx1_p & v85628f;
assign v8558d9 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a31ed;
assign v8a33be = EMPTY_p & v8a3329 | !EMPTY_p & v856992;
assign v844fb1 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & !v844f91;
assign v85be78 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v873899;
assign v8a2e46 = stateG12_p & v8559ee | !stateG12_p & !v844f91;
assign v8a2ae0 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8962c7;
assign v8579da = jx1_p & v8a3183 | !jx1_p & v8a2fba;
assign v8a2837 = ENQ_p & v85741f | !ENQ_p & v85aac2;
assign v855ea7 = EMPTY_p & v856063 | !EMPTY_p & v8a28af;
assign v8557b0 = ENQ_p & v856c57 | !ENQ_p & v85525c;
assign v85605e = jx0_p & v8a2e42 | !jx0_p & !v8a24a6;
assign v855e66 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v876d51;
assign v85eda6 = BtoS_ACK3_p & v844fa0 | !BtoS_ACK3_p & !v844f91;
assign v8738ae = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v856e0b;
assign v8a3116 = BtoS_ACK1_p & v856639 | !BtoS_ACK1_p & v854edf;
assign v8a282b = ENQ_p & v844fa9 | !ENQ_p & !v8a3002;
assign v8a331c = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a314b;
assign v8579f9 = jx1_p & v8a31f6 | !jx1_p & v8574ba;
assign v854151 = jx0_p & v88ac2c | !jx0_p & v856af6;
assign v85edeb = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v85eb9f;
assign v856991 = stateG7_1_p & v855700 | !stateG7_1_p & v856144;
assign v856801 = jx1_p & v85698e | !jx1_p & !v8a31d1;
assign v854fd3 = StoB_REQ0_p & v8a30b3 | !StoB_REQ0_p & !v844f91;
assign v855e36 = jx1_p & v85606a | !jx1_p & !v844f91;
assign v856e4a = ENQ_p & v85741f | !ENQ_p & v854f04;
assign v855a02 = jx1_p & v855f7c | !jx1_p & v856553;
assign v8a3262 = BtoS_ACK0_p & v844fe7 | !BtoS_ACK0_p & v8a33cf;
assign v8a323b = stateG7_1_p & v8a2cce | !stateG7_1_p & v855acb;
assign v8a2ddc = ENQ_p & v8a313f | !ENQ_p & v854a8f;
assign v854b17 = jx0_p & v89cb27 | !jx0_p & v844f91;
assign v8a332b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3270;
assign v8a2c65 = ENQ_p & v88375a | !ENQ_p & v8a307a;
assign v8562a3 = jx0_p & v8a2f9b | !jx0_p & v844f91;
assign v8541c3 = jx1_p & v844fc1 | !jx1_p & !v8a2fac;
assign v8558a0 = StoB_REQ0_p & v854b33 | !StoB_REQ0_p & v856a09;
assign v8a30cd = RtoB_ACK1_p & v855ebf | !RtoB_ACK1_p & v8a2bb4;
assign v854b6c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a33d9;
assign v8566e1 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v870ea9;
assign v8a3315 = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v8a336c;
assign v8a3332 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v856026;
assign v85ab2f = EMPTY_p & v8553d5 | !EMPTY_p & v8564e4;
assign v8a2b29 = EMPTY_p & v8558d2 | !EMPTY_p & v8557cd;
assign v8a3257 = BtoS_ACK1_p & v87c725 | !BtoS_ACK1_p & v855542;
assign v8738de = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a3035;
assign v8a243e = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v854a71;
assign v8a3181 = jx0_p & v854cad | !jx0_p & v856b69;
assign v8a3290 = BtoS_ACK0_p & v8561e1 | !BtoS_ACK0_p & v856b1f;
assign v89cb27 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v8a3393;
assign v8a3080 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8a312e;
assign v8962fa = DEQ_p & v85798c | !DEQ_p & v8a2f08;
assign v8a314c = RtoB_ACK0_p & v857727 | !RtoB_ACK0_p & v854b0e;
assign v855c80 = ENQ_p & v8a31dc | !ENQ_p & v871174;
assign v8575b3 = StoB_REQ2_p & v883730 | !StoB_REQ2_p & v8a331b;
assign v856cce = jx2_p & v8a31ee | !jx2_p & v844f91;
assign v8561c3 = RtoB_ACK1_p & v8a2d5f | !RtoB_ACK1_p & v855047;
assign v8557f6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3053;
assign v85694d = jx0_p & v89626e | !jx0_p & v8a3275;
assign v857452 = BtoS_ACK2_p & v8a3036 | !BtoS_ACK2_p & v8560f5;
assign v856262 = BtoS_ACK1_p & v856422 | !BtoS_ACK1_p & v854a89;
assign v8a33d3 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8685f8;
assign v871154 = jx0_p & v85ecec | !jx0_p & !v844f91;
assign v85eb80 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v867ef3;
assign v8a3120 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3227;
assign v8a3268 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8552f8;
assign v854edf = StoB_REQ1_p & v8630d3 | !StoB_REQ1_p & v865fb9;
assign v8a324a = jx2_p & v87c743 | !jx2_p & !v855046;
assign v89612f = jx1_p & v856786 | !jx1_p & v857547;
assign v8a30c5 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3336;
assign v855bdb = BtoS_ACK0_p & v8711c0 | !BtoS_ACK0_p & v8a3325;
assign v8a3143 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v856b6b;
assign v855a09 = jx0_p & v857979 | !jx0_p & v85698e;
assign v8a302d = DEQ_p & v8554e5 | !DEQ_p & v856c36;
assign v854188 = StoB_REQ3_p & v8a24df | !StoB_REQ3_p & v844f91;
assign v8a2fa6 = BtoS_ACK0_p & v8a3186 | !BtoS_ACK0_p & v8550b4;
assign v8549fe = jx2_p & v85746e | !jx2_p & !v855674;
assign v8a310a = jx1_p & v8a2fd5 | !jx1_p & v8617f7;
assign v855739 = jx0_p & v8a3237 | !jx0_p & v844f91;
assign v8a33de = BtoS_ACK0_p & v854a11 | !BtoS_ACK0_p & v854edc;
assign v85610f = jx2_p & v86f537 | !jx2_p & v8a2eb6;
assign v8a32d9 = jx1_p & v854b14 | !jx1_p & !v855a66;
assign v85520c = jx1_p & v854194 | !jx1_p & v854eb5;
assign v8a3042 = BtoS_ACK0_p & v8a30f6 | !BtoS_ACK0_p & v8a3282;
assign v8a3173 = EMPTY_p & v8557b0 | !EMPTY_p & !v8a31bc;
assign v855dee = jx0_p & v8a3262 | !jx0_p & !v844f9d;
assign v8a3245 = jx0_p & v855bdb | !jx0_p & v8a311b;
assign v85edf0 = BtoS_ACK0_p & v8711c0 | !BtoS_ACK0_p & v8a31b1;
assign v855d52 = jx0_p & v855a9b | !jx0_p & !v8a336b;
assign v854bcd = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8a3232;
assign v855a66 = jx0_p & v8a3393 | !jx0_p & v844f91;
assign v88abc3 = EMPTY_p & v8a329c | !EMPTY_p & v85ab14;
assign v856945 = stateG7_1_p & v844f91 | !stateG7_1_p & v8a33be;
assign v854cd0 = jx1_p & v844f91 | !jx1_p & v8a283c;
assign v8a3327 = BtoS_ACK0_p & v855eb2 | !BtoS_ACK0_p & v8a327d;
assign v855df1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a306f;
assign v8a3066 = DEQ_p & v8a2ef0 | !DEQ_p & v854a55;
assign v8a3273 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v856bea;
assign v8a31c0 = ENQ_p & v85741f | !ENQ_p & v857583;
assign v8552ac = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8a3386;
assign v896167 = DEQ_p & v8a2ef0 | !DEQ_p & v854ccd;
assign v8a3155 = ENQ_p & v87e83a | !ENQ_p & v8a3405;
assign v856cee = jx0_p & v8a3152 | !jx0_p & !v856786;
assign v857583 = jx2_p & v8a2dfb | !jx2_p & v8579da;
assign v8a2b63 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a302a;
assign v85548d = ENQ_p & v8a31dc | !ENQ_p & v8a2c75;
assign v8a31ca = StoB_REQ2_p & v855ef6 | !StoB_REQ2_p & !v844f91;
assign v8a2824 = jx2_p & v8a3189 | !jx2_p & v856b69;
assign v85416e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3257;
assign v85bce8 = jx0_p & v8552ea | !jx0_p & v8a31b8;
assign v8a2b16 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v867273;
assign v8a33ae = jx1_p & v8a2fd5 | !jx1_p & v8a333b;
assign v8a2b82 = StoB_REQ0_p & v85614f | !StoB_REQ0_p & v855ffb;
assign v855c08 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v8a31f4 = jx1_p & v85617a | !jx1_p & v8573a4;
assign v8a3160 = jx2_p & v8a30b0 | !jx2_p & !v85793b;
assign v8a31ad = jx1_p & v854f8b | !jx1_p & !v855a09;
assign v8a30be = ENQ_p & v855f60 | !ENQ_p & v85690e;
assign v854cc4 = jx0_p & v8566c4 | !jx0_p & v8a2fd5;
assign v88b742 = BtoS_ACK2_p & v8a33c1 | !BtoS_ACK2_p & v8a3318;
assign v8a3399 = jx0_p & v8a31d9 | !jx0_p & !v8552c6;
assign v8a338f = jx2_p & v860488 | !jx2_p & !v856d52;
assign v855c02 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v854ee4;
assign v8a3135 = BtoS_ACK2_p & v8567ec | !BtoS_ACK2_p & v8a3166;
assign v8a3079 = ENQ_p & v844fa9 | !ENQ_p & !v855de8;
assign v856df4 = jx0_p & v856c4f | !jx0_p & !v8554aa;
assign v8560ff = jx1_p & v844f91 | !jx1_p & !v8a32b3;
assign v8a3251 = EMPTY_p & v8a31ae | !EMPTY_p & v8551ba;
assign v855065 = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v8552c8;
assign v8a31a7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8555ef;
assign v85555f = EMPTY_p & v855e0f | !EMPTY_p & !v8a2891;
assign v855f5b = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844fad;
assign v8a2e43 = jx2_p & v8a3210 | !jx2_p & v8a2cbd;
assign v8a3265 = StoB_REQ2_p & v8a29a5 | !StoB_REQ2_p & v844f91;
assign v85543e = BtoS_ACK0_p & v8a333a | !BtoS_ACK0_p & v855eb3;
assign v8a30bb = jx1_p & v85606a | !jx1_p & !v855e40;
assign v85509e = jx0_p & v8a3391 | !jx0_p & !v870eb8;
assign v87c729 = jx2_p & v8a323e | !jx2_p & v856047;
assign v8a288c = stateG7_1_p & v8a331a | !stateG7_1_p & v86a9e8;
assign v8a3221 = ENQ_p & v87c729 | !ENQ_p & v856a98;
assign v8563ed = stateG12_p & v85741f | !stateG12_p & v8a2fba;
assign v8569b3 = EMPTY_p & v855b24 | !EMPTY_p & v8a3239;
assign v8551c8 = StoB_REQ1_p & v8a3130 | !StoB_REQ1_p & v85aad7;
assign v88ab9d = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8a31f3;
assign v857a7a = EMPTY_p & v856253 | !EMPTY_p & v88abd1;
assign v8541e8 = jx0_p & v85663b | !jx0_p & v844f9d;
assign v8a2fce = RtoB_ACK0_p & v857414 | !RtoB_ACK0_p & v856b13;
assign v8550a1 = BtoS_ACK0_p & v8a336d | !BtoS_ACK0_p & v896162;
assign v883c9a = ENQ_p & v856b26 | !ENQ_p & v8a2824;
assign v8a2479 = jx0_p & v8a2a05 | !jx0_p & v844f91;
assign v854d35 = BtoS_ACK1_p & v8562d8 | !BtoS_ACK1_p & v8a3356;
assign v8a328a = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v856c01;
assign v8a3236 = DEQ_p & v844f91 | !DEQ_p & v8a32e8;
assign v8a32fb = DEQ_p & v856901 | !DEQ_p & v8617d4;
assign v8a2bfd = jx1_p & v8559f8 | !jx1_p & v876d53;
assign v855016 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v854a89;
assign v8a303b = StoB_REQ1_p & v85ed6f | !StoB_REQ1_p & v855eb2;
assign v8a339f = ENQ_p & v8574ba | !ENQ_p & v8a327f;
assign v8567aa = DEQ_p & v856828 | !DEQ_p & v876d41;
assign v8a32ea = StoB_REQ1_p & v8a29d7 | !StoB_REQ1_p & v854b71;
assign v8a2486 = DEQ_p & v85786a | !DEQ_p & v855f55;
assign v8a30b1 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a0e17;
assign v8a3094 = jx0_p & v8a338c | !jx0_p & v85606a;
assign v855542 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v856500;
assign v883cb2 = BtoS_ACK1_p & v86c421 | !BtoS_ACK1_p & v86c9ca;
assign v8a334e = StoB_REQ1_p & v8a322d | !StoB_REQ1_p & v85ed30;
assign v856007 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a2f6b;
assign v857731 = StoB_REQ4_p & v8a2f21 | !StoB_REQ4_p & v844f91;
assign v8a3090 = jx1_p & v854151 | !jx1_p & v8a3094;
assign v8a31ff = BtoS_ACK2_p & v8a3036 | !BtoS_ACK2_p & v8a316b;
assign v8a2f07 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a3363;
assign v8a336c = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & !v844f9f;
assign v857572 = EMPTY_p & v8a3333 | !EMPTY_p & v855137;
assign v8a312e = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v8685f8;
assign v8a30fc = EMPTY_p & v8a2cc7 | !EMPTY_p & v8a31bb;
assign v8a3053 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a2958;
assign v8a30ab = RtoB_ACK1_p & v8a2898 | !RtoB_ACK1_p & v8a319e;
assign v8a0de5 = stateG7_1_p & v8a28de | !stateG7_1_p & v854a23;
assign v88373a = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v856c9f;
assign v8a3150 = jx0_p & v8a30e7 | !jx0_p & !v844f91;
assign v8a3386 = StoB_REQ1_p & v8555ef | !StoB_REQ1_p & !v844f91;
assign v8a304b = jx1_p & v844f91 | !jx1_p & v8a30fb;
assign v8a2ff2 = FULL_p & v8a339f | !FULL_p & v855fab;
assign v883709 = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v8a31b9;
assign v89614f = EMPTY_p & v8558d2 | !EMPTY_p & v8a3182;
assign v8551dd = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v85ed6f;
assign v85778c = jx1_p & v844f91 | !jx1_p & !v855acd;
assign v8568b1 = StoB_REQ1_p & v87d020 | !StoB_REQ1_p & v861784;
assign v8a31ee = jx1_p & v844f91 | !jx1_p & !v8a33c6;
assign v8774cb = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8549db;
assign v85aab4 = ENQ_p & v85413e | !ENQ_p & v8565c6;
assign v8a3322 = BtoS_ACK1_p & v8a3032 | !BtoS_ACK1_p & v8a29eb;
assign v8a3058 = ENQ_p & v8a3211 | !ENQ_p & v89624b;
assign v8564c9 = StoB_REQ2_p & v85791e | !StoB_REQ2_p & v855114;
assign v857469 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8a31bd;
assign v8a313d = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v85687a;
assign v85ab44 = DEQ_p & v8551f9 | !DEQ_p & v8a336e;
assign v8a3026 = ENQ_p & v844f91 | !ENQ_p & v8a33b0;
assign v8553e6 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a3130;
assign v857b65 = jx0_p & v8a311e | !jx0_p & !v85edeb;
assign v85528e = BtoS_ACK0_p & v88ab81 | !BtoS_ACK0_p & v8a29c6;
assign v8a31c6 = DEQ_p & v896289 | !DEQ_p & v8a315c;
assign v855e1c = BtoS_ACK2_p & v8711d9 | !BtoS_ACK2_p & v85ed6f;
assign v8a31b9 = StoB_REQ1_p & v8a3377 | !StoB_REQ1_p & v8a3096;
assign v855fab = ENQ_p & v8574ba | !ENQ_p & v855b2b;
assign v857aed = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v8a334e;
assign v8a3381 = jx1_p & v856903 | !jx1_p & !v844f91;
assign v856047 = jx1_p & v8a2bd1 | !jx1_p & v8a31d5;
assign v85699f = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v860093;
assign v883733 = jx0_p & v8a330f | !jx0_p & v844f91;
assign v85524b = stateG12_p & v85606a | !stateG12_p & v856786;
assign v8576c3 = EMPTY_p & v8a2f17 | !EMPTY_p & v8a3044;
assign v8a3171 = RtoB_ACK1_p & v8a3117 | !RtoB_ACK1_p & v8a2b29;
assign BtoS_ACK4_n = !v87c76f;
assign v85e12c = BtoR_REQ1_p & v8574ef | !BtoR_REQ1_p & v8a3223;
assign v85a4b4 = DEQ_p & v8a2894 | !DEQ_p & v8a3048;
assign v855d44 = ENQ_p & v856553 | !ENQ_p & !v8a2c53;
assign v8a30aa = jx2_p & v8a304b | !jx2_p & v844f91;
assign v852505 = BtoS_ACK0_p & v844fa0 | !BtoS_ACK0_p & v871675;
assign v870ea7 = jx2_p & v8a329e | !jx2_p & v856624;
assign BtoR_REQ1_n = !v883ce3;
assign v877670 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a29e3;
assign v8a30ba = jx0_p & v854feb | !jx0_p & v844f91;
assign v8a2a8c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v85540d;
assign v856c36 = ENQ_p & v86b41a | !ENQ_p & v867269;
assign v855b2b = jx2_p & v8a3070 | !jx2_p & !v8a3200;
assign v855e45 = stateG12_p & v844fa9 | !stateG12_p & !v844f91;
assign v8a3278 = jx0_p & v8a32b9 | !jx0_p & v844f91;
assign v854eb5 = jx0_p & v856bd6 | !jx0_p & v8550fb;
assign v8a2e76 = RtoB_ACK0_p & v8a24b8 | !RtoB_ACK0_p & v8a320e;
assign v866887 = BtoR_REQ0_p & v8a314c | !BtoR_REQ0_p & v8a2e1f;
assign v883710 = StoB_REQ2_p & v8a0e03 | !StoB_REQ2_p & v85523e;
assign v8a29c6 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a332e;
assign v8579f4 = ENQ_p & v85570e | !ENQ_p & v857583;
assign v856023 = jx0_p & v85ecec | !jx0_p & v85698e;
assign BtoS_ACK2_n = !v8a0e69;
assign v855edc = jx1_p & v8a2c50 | !jx1_p & !v85adee;
assign v85687a = StoB_REQ1_p & v8a318e | !StoB_REQ1_p & v856df1;
assign v85be86 = EMPTY_p & v8a24d1 | !EMPTY_p & !v854994;
assign v844f9d = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v844f91;
assign v8a302f = jx2_p & v8a326d | !jx2_p & v87c763;
assign v8a2e1f = BtoR_REQ1_p & v8550db | !BtoR_REQ1_p & v85be86;
assign v8a31c8 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8555ef;
assign v8a3082 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8560ea;
assign v857917 = StoB_REQ2_p & v85509b | !StoB_REQ2_p & v854f97;
assign v85d4ae = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8a30b1;
assign v85698c = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v8a3077;
assign v8a322c = RtoB_ACK1_p & v856d80 | !RtoB_ACK1_p & v8a32e2;
assign v8a2fc5 = stateG7_1_p & v8a3251 | !stateG7_1_p & v8a3364;
assign v88371a = jx2_p & v856497 | !jx2_p & !v8a2bfd;
assign v8a3050 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8a3360;
assign v8a31ae = ENQ_p & v87c729 | !ENQ_p & v8a2c75;
assign v856e3f = jx1_p & v8a3284 | !jx1_p & v854cc4;
assign v8556c9 = BtoS_ACK0_p & v8711cf | !BtoS_ACK0_p & v855708;
assign v878154 = jx2_p & v8a3134 | !jx2_p & !v8a32d9;
assign v8a312b = BtoS_ACK0_p & v857a31 | !BtoS_ACK0_p & v8552de;
assign v854a07 = DEQ_p & v855fb0 | !DEQ_p & v8a329c;
assign v856372 = EMPTY_p & v855ead | !EMPTY_p & v855a6a;
assign v85562c = DEQ_p & v8a30a6 | !DEQ_p & v856432;
assign v855a4d = RtoB_ACK0_p & v8a32d0 | !RtoB_ACK0_p & v8a0de5;
assign v8a3023 = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v85628e;
assign v8555a0 = jx1_p & v855865 | !jx1_p & !v86624f;
assign v8553e7 = StoB_REQ3_p & v8a2f21 | !StoB_REQ3_p & v85523e;
assign v854a23 = EMPTY_p & v876d41 | !EMPTY_p & v85edc8;
assign v89fce5 = BtoS_ACK0_p & v8a337f | !BtoS_ACK0_p & v8561e7;
assign v856e47 = jx0_p & v8a2ec1 | !jx0_p & v856624;
assign v855e0f = ENQ_p & v87e83a | !ENQ_p & v85525c;
assign v856556 = jx0_p & v89cb27 | !jx0_p & !v870eb8;
assign v8a32f4 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v855311;
assign v85628e = StoB_REQ2_p & v883730 | !StoB_REQ2_p & v856c80;
assign v86dd6d = FULL_p & v876d41 | !FULL_p & v8a2c6e;
assign v8a3346 = RtoB_ACK1_p & v85ab2f | !RtoB_ACK1_p & v8565ef;
assign v856ab3 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v86c421;
assign v8a2b44 = jx2_p & v85ec27 | !jx2_p & v856b69;
assign v85618d = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v85540d;
assign v8a3182 = DEQ_p & v85743a | !DEQ_p & v8a308f;
assign v8a31ab = jx0_p & v8557a6 | !jx0_p & !v85577c;
assign v8a315b = StoB_REQ0_p & v8565de | !StoB_REQ0_p & v844f91;
assign v85ab2e = BtoS_ACK2_p & v856422 | !BtoS_ACK2_p & v8541c6;
assign v87d033 = BtoS_ACK1_p & v8a333a | !BtoS_ACK1_p & v8a32d3;
assign v8a320f = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v8a337d;
assign v855865 = jx0_p & v8558e6 | !jx0_p & !v8a31c5;
assign v854b24 = EMPTY_p & v8568be | !EMPTY_p & v8a30c4;
assign v8556bc = jx1_p & v855e45 | !jx1_p & v844fa9;
assign v8a295f = FULL_p & v855002 | !FULL_p & v8a2a85;
assign v857692 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v8a3081;
assign v8a30ce = jx1_p & v8a331e | !jx1_p & !v856786;
assign v8a31a8 = ENQ_p & v855254 | !ENQ_p & v85576d;
assign v8a3044 = DEQ_p & v85a137 | !DEQ_p & v8a330a;
assign v8554e5 = ENQ_p & v856b26 | !ENQ_p & v8a30f0;
assign v854cf3 = DEQ_p & v8a31af | !DEQ_p & v8a3083;
assign v8a3035 = StoB_REQ0_p & v8a2893 | !StoB_REQ0_p & v844f91;
assign v8554aa = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8a3338;
assign v8a287d = StoB_REQ1_p & v8a32a1 | !StoB_REQ1_p & v844f91;
assign v85ab38 = EMPTY_p & v8a2984 | !EMPTY_p & v855a6a;
assign v8a30fb = jx0_p & v8a30e9 | !jx0_p & !v844f9d;
assign v8a29eb = StoB_REQ1_p & v8a29d7 | !StoB_REQ1_p & !v8a30b8;
assign v89fcfa = jx1_p & v8559f8 | !jx1_p & v844f91;
assign v8a32b3 = jx0_p & v8549e9 | !jx0_p & !v8554aa;
assign v8564e4 = DEQ_p & v85743a | !DEQ_p & v8a296b;
assign v8578b4 = jx1_p & v85ed68 | !jx1_p & !v844f91;
assign v8a3387 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v856651;
assign v8630d3 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856acb;
assign v8573ee = StoB_REQ4_p & v8a2f21 | !StoB_REQ4_p & v844f9f;
assign v8a30c1 = jx1_p & v8a3151 | !jx1_p & v8a300d;
assign v855ddf = jx1_p & v8554f7 | !jx1_p & v856553;
assign v855780 = StoB_REQ0_p & v8a2b19 | !StoB_REQ0_p & v8a30e5;
assign v8962c7 = StoB_REQ2_p & v871051 | !StoB_REQ2_p & v8552b4;
assign v856270 = jx1_p & v855d45 | !jx1_p & v855398;
assign v8a24a6 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8553cf;
assign v8a31dd = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v8a31fe;
assign v8549db = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856e2b;
assign v854c5b = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v854f90;
assign v856901 = ENQ_p & v854b5e | !ENQ_p & v844f91;
assign v8564e9 = ENQ_p & v85413e | !ENQ_p & v8a2824;
assign v8703da = jx1_p & v856903 | !jx1_p & v871154;
assign v856438 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8a2c94;
assign v8a331b = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v85635c;
assign v857b42 = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v8a32af;
assign v8617f7 = jx0_p & v856966 | !jx0_p & v8a3273;
assign v8a3234 = DEQ_p & v8554e5 | !DEQ_p & v856432;
assign v8558d2 = ENQ_p & v844f91 | !ENQ_p & !v855658;
assign v8a33c0 = jx2_p & v8a30c1 | !jx2_p & v855df9;
assign v8557cd = DEQ_p & v85743a | !DEQ_p & v8a3088;
assign v857aee = jx1_p & v85606a | !jx1_p & !v8567ad;
assign v855e5a = RtoB_ACK1_p & v86aa1f | !RtoB_ACK1_p & v85a3a3;
assign v8554d7 = EMPTY_p & v8a30af | !EMPTY_p & v8a3234;
assign v896174 = RtoB_ACK0_p & v855ce1 | !RtoB_ACK0_p & v87c747;
assign v8a33c2 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v86aa4b;
assign v869f3f = StoB_REQ1_p & v8a3314 | !StoB_REQ1_p & v8a319c;
assign v8541e6 = jx0_p & v8a2fb0 | !jx0_p & v854fa7;
assign v8a28de = RtoB_ACK1_p & v8a32d0 | !RtoB_ACK1_p & v854a23;
assign v857a8c = ENQ_p & v844f91 | !ENQ_p & !v8a33c0;
assign v8a331f = ENQ_p & v855298 | !ENQ_p & v870ea7;
assign v856063 = ENQ_p & v855254 | !ENQ_p & v844f91;
assign v8962e0 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v88372d;
assign v8a3249 = BtoS_ACK0_p & v857880 | !BtoS_ACK0_p & v8a2dc2;
assign v8711c0 = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v8a3086;
assign v854b0e = stateG7_1_p & v87c6f7 | !stateG7_1_p & v8a32d7;
assign v8a323a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v857619;
assign v8a30e2 = jx1_p & v8a31b2 | !jx1_p & v856556;
assign v85aac2 = jx2_p & v8a3108 | !jx2_p & v8565a7;
assign v854feb = BtoS_ACK0_p & v855c79 | !BtoS_ACK0_p & v86938f;
assign v854aa0 = jx2_p & v858911 | !jx2_p & v8711ac;
assign v85413d = BtoS_ACK0_p & v8a3129 | !BtoS_ACK0_p & v896106;
assign v8559f8 = jx0_p & v8a311e | !jx0_p & v844f91;
assign v8a2f46 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v873fa6;
assign v86a9c5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a338c;
assign v855a2a = stateG12_p & v844fa9 | !stateG12_p & !v8a2fd5;
assign v872af1 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v8711d9;
assign v86180e = BtoR_REQ0_p & v86a9dc | !BtoR_REQ0_p & v85679c;
assign v8962f6 = DEQ_p & v896289 | !DEQ_p & v855002;
assign v8549e9 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v855147;
assign v8a310d = ENQ_p & v8574eb | !ENQ_p & v8a2bb0;
assign v8a3305 = StoB_REQ0_p & v8556d0 | !StoB_REQ0_p & v844f91;
assign v8a3292 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8a3241;
assign v8a332c = jx1_p & v85ed68 | !jx1_p & v883725;
assign v855845 = EMPTY_p & v854a55 | !EMPTY_p & v8a30e1;
assign v8a3307 = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v856df1;
assign v856af6 = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v8a32f8;
assign v876d53 = jx0_p & v8a0e4f | !jx0_p & !v844f91;
assign v8a337d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854a53;
assign v86a9f3 = StoB_REQ0_p & v85eb80 | !StoB_REQ0_p & v844f91;
assign v8a33d8 = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v8a332b;
assign v8a3237 = BtoS_ACK0_p & v8a3379 | !BtoS_ACK0_p & v86c364;
assign v8a3089 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v8a3355 = BtoS_ACK0_p & v855311 | !BtoS_ACK0_p & v857651;
assign v85edc8 = DEQ_p & v866b88 | !DEQ_p & v876d41;
assign v8a29d0 = jx1_p & v854194 | !jx1_p & v86550e;
assign v854b5f = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a331b;
assign v8a33ad = jx0_p & v856653 | !jx0_p & !v854194;
assign v85795e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8552ac;
assign v8a316b = StoB_REQ2_p & v856e2b | !StoB_REQ2_p & v854c40;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v89629f = BtoS_ACK2_p & v88b745 | !BtoS_ACK2_p & v856731;
assign v8a3263 = jx1_p & v85698e | !jx1_p & !v8a3392;
assign v8a31e2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v85576e;
assign v8a31d2 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v883cad;
assign v8560a3 = RtoB_ACK1_p & v855bec | !RtoB_ACK1_p & v875b8c;
assign v8a3219 = jx0_p & v8a30e9 | !jx0_p & !v8a3159;
assign v8a2fb0 = BtoS_ACK0_p & v8a336d | !BtoS_ACK0_p & v8a304e;
assign v87c759 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v8a31c8;
assign v8a32c6 = ENQ_p & v844fa9 | !ENQ_p & !v8a3244;
assign v85522b = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3025;
assign v876345 = jx2_p & v873280 | !jx2_p & !v857624;
assign v8568be = ENQ_p & v844f91 | !ENQ_p & !v8a31c7;
assign v85d533 = jx0_p & v8558cf | !jx0_p & v8a32a3;
assign v8a31b2 = jx0_p & v857b70 | !jx0_p & !v8a31e4;
assign v871051 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8a3315;
assign v8a24d1 = ENQ_p & v856c57 | !ENQ_p & v878154;
assign v8a3363 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8a33d3;
assign v8a2e8b = jx1_p & v844f91 | !jx1_p & v8a2d89;
assign v8a329e = jx1_p & v844f91 | !jx1_p & !v8a3372;
assign v8575a5 = jx2_p & v8a30b7 | !jx2_p & v855386;
assign v8a2eb6 = jx1_p & v8a3043 | !jx1_p & v844f91;
assign v86179a = EMPTY_p & v8a31c0 | !EMPTY_p & v8575fe;
assign v89625f = BtoS_ACK3_p & v855b05 | !BtoS_ACK3_p & v8a33c1;
assign v8575fe = DEQ_p & v8579f4 | !DEQ_p & v854ccd;
assign v854ed3 = StoB_REQ2_p & v8a308c | !StoB_REQ2_p & !v872af1;
assign v856ad7 = StoB_REQ1_p & v8a32c4 | !StoB_REQ1_p & v844f91;
assign v8a3288 = RtoB_ACK0_p & v854fe9 | !RtoB_ACK0_p & v8a323b;
assign v8553de = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v854ef2;
assign v8552b8 = StoB_REQ0_p & v8573cd | !StoB_REQ0_p & v8a309a;
assign v8a2c53 = jx2_p & v855ebc | !jx2_p & !v8a31ad;
assign v854fa7 = BtoS_ACK0_p & v8564d2 | !BtoS_ACK0_p & v8a3362;
assign v857969 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a333a;
assign v8a3285 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86aa49;
assign v86a9cf = jx2_p & v8836fc | !jx2_p & !v8a30ce;
assign v86fe32 = jx2_p & v854a06 | !jx2_p & v856624;
assign v855060 = ENQ_p & v8a332a | !ENQ_p & !v8574e2;
assign v8a33db = jx0_p & v8a3250 | !jx0_p & v844f91;
assign v85419c = jx0_p & v8a3393 | !jx0_p & !v870eb8;
assign v8a332a = jx2_p & v855a02 | !jx2_p & v856553;
assign v8a30b7 = jx1_p & v8a3151 | !jx1_p & v87532a;
assign v8a31dc = jx2_p & v8a30bb | !jx2_p & v856047;
assign v854ef2 = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v856c23;
assign v873756 = RtoB_ACK1_p & v857b51 | !RtoB_ACK1_p & v855998;
assign v8a3153 = jx0_p & v8a3250 | !jx0_p & !v8a24a6;
assign v8a311b = BtoS_ACK0_p & v85ed6f | !BtoS_ACK0_p & v8a31cc;
assign v8a2fac = jx0_p & v8a29ad | !jx0_p & v844f91;
assign v8a31bb = DEQ_p & v855060 | !DEQ_p & v8a295f;
assign v8565c6 = jx2_p & v854c44 | !jx2_p & v87c763;
assign v8559ce = BtoS_ACK1_p & v854a11 | !BtoS_ACK1_p & v8557be;
assign v856781 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85e22c;
assign v85648f = RtoB_ACK0_p & v8a2be7 | !RtoB_ACK0_p & !v8a32fe;
assign v8a3196 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v86a9f3;
assign v8551a3 = jx0_p & v85663b | !jx0_p & v8a311b;
assign v857979 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8a30b3;
assign v8a2d10 = jx1_p & v844fc1 | !jx1_p & v8a311d;
assign v87116a = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v854a0a;
assign v856790 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v854c76;
assign v854a55 = ENQ_p & v85741f | !ENQ_p & v844f91;
assign v857b51 = EMPTY_p & v8a326c | !EMPTY_p & v8556ec;
assign v85ab2a = StoB_REQ1_p & v85754a | !StoB_REQ1_p & v855564;
assign v85698e = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8552e8;
assign v8a3186 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v8552e8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a30b3;
assign v88ab81 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v8a2daf = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v857a54;
assign v857a4d = jx0_p & v8a3262 | !jx0_p & !v8a3159;
assign v855492 = jx0_p & v857932 | !jx0_p & v856441;
assign v8a32fe = stateG7_1_p & v844fa3 | !stateG7_1_p & !v844f91;
assign v855790 = StoB_REQ3_p & v8a2f21 | !StoB_REQ3_p & v857731;
assign v8a302a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v856be3;
assign v855c6b = BtoS_ACK1_p & v8a333a | !BtoS_ACK1_p & v857534;
assign v8a296b = FULL_p & v844f91 | !FULL_p & v8a32e8;
assign v86c425 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v8551d0;
assign v8560c5 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & !v86c425;
assign v883741 = ENQ_p & v856aa1 | !ENQ_p & v8a2e43;
assign v856acb = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a2f21;
assign v855ed8 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8565b9;
assign v8a3140 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a2935;
assign v8a32e2 = EMPTY_p & v88ab43 | !EMPTY_p & v855182;
assign v854aed = RtoB_ACK1_p & v855db2 | !RtoB_ACK1_p & v844f91;
assign v857aaa = ENQ_p & v85413e | !ENQ_p & v883cb8;
assign v8a311d = jx0_p & v8a3045 | !jx0_p & v8a3235;
assign v856e2b = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v854bf7;
assign v856253 = ENQ_p & v85413e | !ENQ_p & v857783;
assign v8a304d = jx1_p & v883733 | !jx1_p & !v88ab84;
assign v856828 = ENQ_p & v8a302e | !ENQ_p & !v8566b8;
assign v85554c = BtoR_REQ1_p & v8a2fce | !BtoR_REQ1_p & v856c8d;
assign v856883 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a337f;
assign v855565 = stateG12_p & v85413e | !stateG12_p & v844f91;
assign v8a32c4 = BtoS_ACK2_p & v88b745 | !BtoS_ACK2_p & v8a302a;
assign v8a3110 = DEQ_p & v856828 | !DEQ_p & v8a335a;
assign v855ffb = BtoS_ACK1_p & v8a3170 | !BtoS_ACK1_p & v88abdb;
assign v855e06 = ENQ_p & v8a313f | !ENQ_p & v8a32b8;
assign v8a309e = EMPTY_p & v8a28c6 | !EMPTY_p & v8a3197;
assign v875b8c = EMPTY_p & v856e4a | !EMPTY_p & v8575fe;
assign v8a2e4a = StoB_REQ2_p & v860093 | !StoB_REQ2_p & v8a304f;
assign v855a9b = BtoS_ACK0_p & v8a3379 | !BtoS_ACK0_p & v8558a0;
assign v8a3164 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8560aa;
assign v8a32ce = jx2_p & v857543 | !jx2_p & v8a31f2;
assign v870d30 = jx1_p & v8a315e | !jx1_p & v85575f;
assign v8a2e89 = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v8a28b9;
assign v8a308c = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f9d;
assign v8a328e = RtoB_ACK0_p & v8a2fc5 | !RtoB_ACK0_p & v856991;
assign v870eba = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v857917;
assign v856195 = jx1_p & v844f91 | !jx1_p & v8a3415;
assign v8a329f = jx2_p & v8a334f | !jx2_p & !v8a317f;
assign v855046 = jx1_p & v855bc8 | !jx1_p & !v85a071;
assign v8a3347 = jx1_p & v85698e | !jx1_p & !v8541e6;
assign v856500 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v868e49;
assign v87c743 = jx1_p & v844f91 | !jx1_p & !v856288;
assign v8566c4 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v854fd3;
assign v854e79 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & !v844f91;
assign v8565a7 = jx1_p & v8a314d | !jx1_p & v856374;
assign v8a30fd = BtoS_ACK2_p & v8567ec | !BtoS_ACK2_p & v883710;
assign v8a2d94 = jx1_p & v855426 | !jx1_p & !v8a334a;
assign v855182 = DEQ_p & v8a3038 | !DEQ_p & v855850;
assign v8562f8 = BtoS_ACK0_p & v8a336d | !BtoS_ACK0_p & v856197;
assign v855001 = jx1_p & v857b65 | !jx1_p & !v8961ce;
assign v854fe9 = EMPTY_p & v8569fe | !EMPTY_p & v85678b;
assign v883cad = BtoS_ACK1_p & v8a337f | !BtoS_ACK1_p & v8a3332;
assign v8575b5 = jx2_p & v8a3398 | !jx2_p & v8a326b;
assign v87c300 = jx1_p & v844f91 | !jx1_p & !v85605e;
assign v8a28c6 = ENQ_p & v855298 | !ENQ_p & v8a32ce;
assign v871174 = jx2_p & v856003 | !jx2_p & v8a3090;
assign v88b745 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844f9d;
assign v85798c = ENQ_p & v857a8e | !ENQ_p & v855e7a;
assign v8a31b6 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v89629f;
assign v8a2dfa = stateG12_p & v85413e | !stateG12_p & v856b69;
assign v876a61 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854ae5;
assign v8a338b = StoB_REQ0_p & v8565b9 | !StoB_REQ0_p & v854ba4;
assign v857b70 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8a3163;
assign v856e7b = StoB_REQ0_p & v854b1a | !StoB_REQ0_p & v8579a9;
assign v8a2d5f = EMPTY_p & v855ead | !EMPTY_p & v855cfe;
assign v8a3184 = StoB_REQ2_p & v8a2c6b | !StoB_REQ2_p & v872af1;
assign v8555b7 = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v88a458;
assign v855a7a = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a0e03;
assign v8a326f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8a31dd;
assign v8a3025 = BtoS_ACK1_p & v87c725 | !BtoS_ACK1_p & v856871;
assign v8565ef = EMPTY_p & v8553d5 | !EMPTY_p & v8557cd;
assign v8a337e = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8541c6;
assign v856ab0 = stateG7_1_p & v8a33bc | !stateG7_1_p & v85a3c4;
assign v856003 = jx1_p & v85606a | !jx1_p & !v85d533;
assign v8a32a1 = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v8a3287;
assign v8a3038 = ENQ_p & v8565ba | !ENQ_p & v8a2bb0;
assign v8a30d5 = EMPTY_p & v8a2cc7 | !EMPTY_p & v855cc1;
assign v857785 = BtoS_ACK2_p & v856422 | !BtoS_ACK2_p & !v856710;
assign v85617a = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8552b8;
assign v8a31cb = stateG7_1_p & v873866 | !stateG7_1_p & v88ab9b;
assign v8a32a7 = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v8573b7;
assign v867273 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v8a2c6b;
assign v8a3074 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v873869;
assign v855cc1 = DEQ_p & v855060 | !DEQ_p & v8a315c;
assign v8a3098 = BtoS_ACK0_p & v8a3129 | !BtoS_ACK0_p & v857ad0;
assign v873613 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a324c;
assign v855de8 = jx2_p & v8a3091 | !jx2_p & v856e3f;
assign v8a33b3 = StoB_REQ2_p & v8a3082 | !StoB_REQ2_p & v856041;
assign v8a2c50 = jx0_p & v856aac | !jx0_p & !v8a30c7;
assign v88ab99 = stateG7_1_p & v8a2d12 | !stateG7_1_p & v8a3016;
assign v855c77 = jx1_p & v856b69 | !jx1_p & v855dee;
assign v8541c6 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8a32ba;
assign v86550e = jx0_p & v8578fc | !jx0_p & v8550fb;
assign v8a33b2 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & !v85635c;
assign v856b69 = BtoS_ACK0_p & v856883 | !BtoS_ACK0_p & v8561e7;
assign v88ab84 = jx0_p & v8a3391 | !jx0_p & v844f91;
assign v855f7c = stateG12_p & v856553 | !stateG12_p & !v85698e;
assign v8a3101 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a2aed;
assign v856c4f = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8a2fe8;
assign v844faf = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v855f60 = jx2_p & v855e36 | !jx2_p & v844f91;
assign v8a2958 = StoB_REQ1_p & v89629f | !StoB_REQ1_p & v844f91;
assign v8a2b42 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a323a;
assign v8a2a91 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v8a3107;
assign v86aa1f = EMPTY_p & v856432 | !EMPTY_p & v8a3198;
assign v855af2 = DEQ_p & v844f91 | !DEQ_p & v85640f;
assign v8a3340 = StoB_REQ0_p & v8a31a7 | !StoB_REQ0_p & !v8a3074;
assign v87c707 = ENQ_p & v8574ba | !ENQ_p & v855935;
assign v8a0e4e = EMPTY_p & v8a28c6 | !EMPTY_p & v85ab44;
assign v8a312d = RtoB_ACK0_p & v8662d9 | !RtoB_ACK0_p & v88ab99;
assign v8a3300 = jx1_p & v8a2fba | !jx1_p & v85694d;
assign v85510d = jx0_p & v8a312b | !jx0_p & !v8a33de;
assign v858bbc = jx2_p & v86f537 | !jx2_p & v89fcfa;
assign v85676f = BtoS_ACK0_p & v856883 | !BtoS_ACK0_p & v855c9e;
assign v8a31df = EMPTY_p & v8a307c | !EMPTY_p & !v8a31bc;
assign v8a32af = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a32a9;
assign v856c23 = BtoS_ACK2_p & v8711d9 | !BtoS_ACK2_p & v8a299a;
assign v8a0e4f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v8a3393;
assign v854f1c = EMPTY_p & v8558fa | !EMPTY_p & v8a3066;
assign v856ad5 = jx1_p & v844f91 | !jx1_p & v8562a3;
assign v8a3232 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v844f91;
assign v855f95 = ENQ_p & v8a324a | !ENQ_p & v8a30d3;
assign v8a2ee2 = jx2_p & v85762e | !jx2_p & !v8a30ce;
assign v8a31e3 = stateG7_1_p & v857595 | !stateG7_1_p & v896294;
assign v8a3227 = StoB_REQ2_p & v855033 | !StoB_REQ2_p & v844f91;
assign v8a30f6 = StoB_REQ1_p & v88ab81 | !StoB_REQ1_p & v8a3032;
assign v8a335a = ENQ_p & v844fa9 | !ENQ_p & !v8a309b;
assign v8560fa = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v855e79;
assign v8556d0 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v86a9eb;
assign v8a333b = jx0_p & v856966 | !jx0_p & v856434;
assign v855cfe = DEQ_p & v8563cf | !DEQ_p & v8541c7;
assign v855ab2 = RtoB_ACK1_p & v8a30fc | !RtoB_ACK1_p & v8a30d5;
assign v856c8d = RtoB_ACK0_p & v88abc3 | !RtoB_ACK0_p & v8a2c62;
assign v8a3294 = ENQ_p & v856553 | !ENQ_p & v8566b6;
assign v8a30b5 = ENQ_p & v86b41a | !ENQ_p & v883cb8;
assign v8a30dc = stateG7_1_p & v8a30f8 | !stateG7_1_p & !v844f91;
assign v89626e = BtoS_ACK0_p & v8a2972 | !BtoS_ACK0_p & v856417;
assign v8a2d89 = jx0_p & v855014 | !jx0_p & !v844f9d;
assign v856624 = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v855eb3;
assign BtoR_REQ0_n = !v8962ff;
assign v8a2891 = DEQ_p & v883741 | !DEQ_p & v855ae0;
assign v85651f = ENQ_p & v85413e | !ENQ_p & v8a30a3;
assign v8566e6 = jx0_p & v855014 | !jx0_p & !v8a3159;
assign v857783 = jx2_p & v8541a9 | !jx2_p & v870d30;
assign v8a315c = FULL_p & v8a329c | !FULL_p & v8a3294;
assign v85613d = BtoS_ACK0_p & v856ab3 | !BtoS_ACK0_p & v8a328b;
assign v8a2984 = ENQ_p & v8574ba | !ENQ_p & v8a321e;
assign v8a2bb4 = EMPTY_p & v8a3079 | !EMPTY_p & v85566d;
assign v85554e = stateG7_1_p & v8a3302 | !stateG7_1_p & v8711bb;
assign v8a2d62 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v883730;
assign v855faf = jx0_p & v8551f8 | !jx0_p & !v8a33d8;
assign v8a24b8 = EMPTY_p & v8a3079 | !EMPTY_p & v8a3110;
assign v85796e = jx0_p & v8a3164 | !jx0_p & v855254;
assign v8a0e55 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v857521;
assign v8560ec = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v854a71;
assign v8a2d78 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v856302;
assign v854b1a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v855a7a;
assign v8a3194 = BtoS_ACK0_p & v856883 | !BtoS_ACK0_p & v856007;
assign v85ed30 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a3128;
assign v8a31d0 = jx2_p & v854cb1 | !jx2_p & v856d52;
assign v8a334a = jx0_p & v8a30e7 | !jx0_p & v8a2fd5;
assign v8549c4 = EMPTY_p & v8a333f | !EMPTY_p & v8a3044;
assign v8a3226 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v855d5e;
assign v856aac = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v85778e;
assign v85508c = jx2_p & v8a31ee | !jx2_p & v856624;
assign v856bfd = RtoB_ACK0_p & v8559bc | !RtoB_ACK0_p & v87116e;
assign v8a326d = jx1_p & v856b69 | !jx1_p & v8a3219;
assign v8a3016 = EMPTY_p & v85579f | !EMPTY_p & v8a3040;
assign v85754a = BtoS_ACK2_p & v8711d9 | !BtoS_ACK2_p & v8a3184;
assign v8a313e = FULL_p & v8a2fd8 | !FULL_p & v865746;
assign v844f9f = StoB_REQ5_p & v844f91 | !StoB_REQ5_p & !v844f91;
assign v856b6b = BtoS_ACK1_p & v8a2972 | !BtoS_ACK1_p & v8a3120;
assign v883725 = jx0_p & v85ecec | !jx0_p & !v8a2fd5;
assign v8a30dd = RtoB_ACK1_p & v855a47 | !RtoB_ACK1_p & v8a3022;
assign v8a327d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a30fe;
assign v855998 = EMPTY_p & v8a326c | !EMPTY_p & v85743c;
assign v8a3106 = stateG12_p & v855254 | !stateG12_p & v844f91;
assign v8a289a = jx1_p & v8563ed | !jx1_p & v85741f;
assign v86f804 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8551d0;
assign v8a3217 = BtoS_ACK3_p & v85523e | !BtoS_ACK3_p & v855790;
assign v855fdf = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v854b7c;
assign v856b8f = FULL_p & v856063 | !FULL_p & v8617d4;
assign v8a321f = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v855c02;
assign v8a3130 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85791e;
assign v8a3317 = jx1_p & v8a2e46 | !jx1_p & v8a311d;
assign v8551f8 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v855780;
assign v856bc0 = StoB_REQ1_p & v8a2d93 | !StoB_REQ1_p & v844f91;
assign v86007c = jx2_p & v8a3263 | !jx2_p & !v855196;
assign v8a3377 = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8a308c;
assign v8573e8 = BtoS_ACK0_p & v8711cf | !BtoS_ACK0_p & v855c3a;
assign v85576d = jx2_p & v855ba9 | !jx2_p & v856270;
assign v8961d4 = BtoR_REQ0_p & v8558ef | !BtoR_REQ0_p & v8a308b;
assign v854b71 = BtoS_ACK2_p & v856422 | !BtoS_ACK2_p & !v8a3334;
assign v8a3054 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v85675f;
assign v8a2cce = RtoB_ACK1_p & v8549ee | !RtoB_ACK1_p & v8569b3;
assign v855398 = jx0_p & v85543e | !jx0_p & v856624;
assign v86a9cb = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v85699f;
assign v8a330f = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v88373a;
assign v8617c9 = DEQ_p & v8a2894 | !DEQ_p & v8541c7;
assign v855879 = BtoS_ACK0_p & v85ed6f | !BtoS_ACK0_p & v876a61;
assign v8a3361 = BtoS_ACK0_p & v8564d2 | !BtoS_ACK0_p & v855397;
assign v8a325f = jx0_p & v85d4ae | !jx0_p & v844f9d;
assign v85509b = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844fb1;
assign v8a2a85 = ENQ_p & v856553 | !ENQ_p & v8a31d0;
assign v8a316d = StoB_REQ1_p & v85698c | !StoB_REQ1_p & v844f91;
assign v854b7c = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v856422;
assign v8560f5 = StoB_REQ2_p & v8a3232 | !StoB_REQ2_p & v854e79;
assign v86aa64 = BtoR_REQ0_p & v855069 | !BtoR_REQ0_p & v856264;
assign v8a3118 = EMPTY_p & v855d44 | !EMPTY_p & v8a31c6;
assign v855bec = EMPTY_p & v856e4a | !EMPTY_p & v854d07;
assign v855386 = jx1_p & v8a31ab | !jx1_p & v8573d3;
assign v855f43 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a321f;
assign v855db2 = EMPTY_p & v844fbd | !EMPTY_p & !v844fbf;
assign v855311 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v844f9b;
assign v856431 = BtoS_ACK0_p & v8a303b | !BtoS_ACK0_p & v8a3301;
assign v855870 = jx0_p & v8a3345 | !jx0_p & v856434;
assign v8a31fb = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v855783;
assign v855f3f = ENQ_p & v855254 | !ENQ_p & v86fe32;
assign v8a3408 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v856349;
assign v863beb = jx1_p & v844f91 | !jx1_p & !v8552f4;
assign v8a3002 = jx2_p & v855d84 | !jx2_p & v8a0dfa;
assign v857487 = ENQ_p & v855298 | !ENQ_p & v855709;
assign v85586d = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3350;
assign v856786 = BtoS_ACK0_p & v855361 | !BtoS_ACK0_p & v856651;
assign v86e908 = stateG7_1_p & v8561c3 | !stateG7_1_p & v86aa4a;
assign v861800 = EMPTY_p & v8a2837 | !EMPTY_p & v896167;
assign v8a3242 = jx0_p & v854feb | !jx0_p & v8573e8;
assign v8a32f8 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v86f804;
assign v8a304f = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v85edc7;
assign v896107 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v88b742;
assign v8a30e7 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a30b3;
assign v8557e1 = jx0_p & v8a3233 | !jx0_p & !v844f9d;
assign v855a89 = BtoS_ACK1_p & v856639 | !BtoS_ACK1_p & v8a2faa;
assign v8a2a3d = StoB_REQ2_p & v856acb | !StoB_REQ2_p & v8559d2;
assign v856c06 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v854b7c;
assign v8a2893 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a318e;
assign v854b2f = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8a2d62;
assign v8a3151 = BtoS_ACK0_p & v855fdf | !BtoS_ACK0_p & !v85531b;
assign v8a3097 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v857785;
assign v8552f4 = jx0_p & v88ab9d | !jx0_p & !v8554aa;
assign v8a2c6c = StoB_REQ1_p & v8a2c94 | !StoB_REQ1_p & !v844f91;
assign v85504a = FULL_p & v8a308f | !FULL_p & v8a3026;
assign v8a2d12 = RtoB_ACK1_p & v8558cb | !RtoB_ACK1_p & v8a28d0;
assign v8a3301 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a306e;
assign v8a31d9 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v85eb80;
assign v8549ee = EMPTY_p & v8a2ddc | !EMPTY_p & v8a2c28;
assign v856636 = StoB_REQ2_p & v856543 | !StoB_REQ2_p & v868e49;
assign v8a31a1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v854a11;
assign v855126 = stateG7_1_p & v8576c3 | !stateG7_1_p & v8549c4;
assign v855ee6 = StoB_REQ3_p & v844fb1 | !StoB_REQ3_p & !v844f91;
assign v855f55 = FULL_p & v8a335a | !FULL_p & v856d91;
assign v8a31e4 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v856176;
assign v85658a = jx2_p & v85659e | !jx2_p & v856d52;
assign v8a299a = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v872af1;
assign v8a2bd1 = jx0_p & v857b42 | !jx0_p & v8a317b;
assign v8a32ae = jx2_p & v8a3380 | !jx2_p & !v8578b4;
assign v856710 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a32ba;
assign v8a3299 = RtoB_ACK0_p & v855c38 | !RtoB_ACK0_p & v8a287f;
assign v87d020 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856790;
assign v86917e = jx1_p & v8a2fba | !jx1_p & v855492;
assign v8a321c = BtoS_ACK1_p & v8a2972 | !BtoS_ACK1_p & v86f89c;
assign v86cbc9 = jx2_p & v873280 | !jx2_p & v844f91;
assign v856b1f = StoB_REQ0_p & v8a2b16 | !StoB_REQ0_p & v8555b7;
assign v8617d4 = ENQ_p & v855254 | !ENQ_p & v856cce;
assign v8a338e = ENQ_p & v8565ba | !ENQ_p & v86a9cf;
assign v85762e = jx1_p & v85606a | !jx1_p & v8541e8;
assign v844fa3 = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v8576bc = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a2cab;
assign v856e00 = BtoS_ACK0_p & v855311 | !BtoS_ACK0_p & v8a32fd;
assign v8a3134 = jx1_p & v844f91 | !jx1_p & v8558d6;
assign v8562af = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855065;
assign v8a3210 = jx1_p & v844fc1 | !jx1_p & !v8a3278;
assign v8574e2 = jx2_p & v8a3347 | !jx2_p & !v856d52;
assign v8550af = stateG7_1_p & v844f91 | !stateG7_1_p & v86f7aa;
assign v855d34 = StoB_REQ2_p & v8a2c6b | !StoB_REQ2_p & v844f91;
assign v896275 = jx0_p & v868cba | !jx0_p & v8a3151;
assign v8a2489 = jx0_p & v8a3042 | !jx0_p & !v8a33cd;
assign v856e74 = EMPTY_p & v8a31a8 | !EMPTY_p & v8a3279;
assign v854e8e = jx1_p & v844f91 | !jx1_p & !v855d52;
assign v856422 = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f9d;
assign v8a3112 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v856438;
assign v854bf7 = BtoS_ACK4_p & v857731 | !BtoS_ACK4_p & v8a2f21;
assign v8a3342 = jx2_p & v88abca | !jx2_p & v85741f;
assign v8a308b = BtoR_REQ1_p & v8557f8 | !BtoR_REQ1_p & v855957;
assign v8a30ef = jx2_p & v85aaf7 | !jx2_p & v8a29f8;
assign v855b2c = jx2_p & v856801 | !jx2_p & !v8a31ad;
assign v88ac2c = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v85eae9;
assign v8a3398 = jx1_p & v844fc1 | !jx1_p & !v85747f;
assign v854cb1 = jx1_p & v844f91 | !jx1_p & v8a31aa;
assign v8a33d9 = BtoS_ACK1_p & v8a2972 | !BtoS_ACK1_p & v854ff9;
assign v8a30bd = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a339a;
assign v8566b8 = jx2_p & v856545 | !jx2_p & v8711ac;
assign v856562 = BtoS_ACK3_p & v844fa0 | !BtoS_ACK3_p & v855b05;
assign v883cb1 = BtoS_ACK1_p & v87c725 | !BtoS_ACK1_p & v8a3408;
assign v8a3326 = EMPTY_p & v855f3f | !EMPTY_p & v8961a7;
assign v86a9eb = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v855033;
assign v8a302c = jx2_p & v8579f9 | !jx2_p & v8574ba;
assign v8a0de9 = BtoS_ACK0_p & v855c08 | !BtoS_ACK0_p & v85795e;
assign v883ce3 = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v856737;
assign v854c44 = jx1_p & v856b69 | !jx1_p & v8566e6;
assign v8836fc = jx1_p & v856786 | !jx1_p & v8550be;
assign v8a2cbd = jx1_p & v856982 | !jx1_p & !v854b17;
assign v8a2e72 = jx1_p & v85565b | !jx1_p & v855254;
assign v856dec = stateG7_1_p & v873853 | !stateG7_1_p & v8a3326;
assign v8a3239 = DEQ_p & v88ab6c | !DEQ_p & v8a330a;
assign v8a3279 = DEQ_p & v8551f9 | !DEQ_p & v856063;
assign v855254 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a2f46;
assign v855cd0 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & v86f804;
assign v856436 = StoB_REQ0_p & v855600 | !StoB_REQ0_p & v8a318a;
assign v8a3250 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8553e6;
assign v8a2dbf = StoB_REQ3_p & v8560ea | !StoB_REQ3_p & !v844f91;
assign v8a3163 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v856648;
assign v8a334f = jx1_p & v844f91 | !jx1_p & !v8563c1;
assign v856966 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v855aec;
assign v8556c1 = jx1_p & v856624 | !jx1_p & !v8a327a;
assign v8a32cc = BtoS_ACK0_p & v855311 | !BtoS_ACK0_p & v896248;
assign v8961cb = RtoB_ACK0_p & v855e27 | !RtoB_ACK0_p & v855126;
assign v8a3027 = EMPTY_p & v8a30cf | !EMPTY_p & !v854fc7;
assign v85531c = EMPTY_p & v8568b8 | !EMPTY_p & !v8a31bc;
assign v89624b = jx2_p & v8a334f | !jx2_p & !v8a332c;
assign v8a31c5 = BtoS_ACK0_p & v856c06 | !BtoS_ACK0_p & v8a3226;
assign v8567ad = jx0_p & v8558cf | !jx0_p & v8556c9;
assign v857ad0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a2d29;
assign v855528 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a31fe;
assign v854d31 = ENQ_p & v856553 | !ENQ_p & !v8574e2;
assign v8a297d = jx1_p & v856cd1 | !jx1_p & !v844f91;
assign v8550e8 = BtoS_ACK0_p & v8a2972 | !BtoS_ACK0_p & v8a3143;
assign v8a30d3 = jx2_p & v8a329b | !jx2_p & !v8a30e2;
assign v8a335b = jx0_p & v8a30eb | !jx0_p & !v844f9d;
assign v8a32ef = RtoB_ACK0_p & v855db2 | !RtoB_ACK0_p & v8a30dc;
assign v85586a = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v8a29dc;
assign v854b8e = BtoS_ACK0_p & v8a31a1 | !BtoS_ACK0_p & v854cbb;
assign v8579c7 = jx0_p & v8550a1 | !jx0_p & v854fa7;
assign v8a30af = ENQ_p & v85413e | !ENQ_p & v8a302f;
assign v854f20 = BtoS_ACK1_p & v87c725 | !BtoS_ACK1_p & v86b201;
assign v854c5c = StoB_REQ2_p & v856790 | !StoB_REQ2_p & v8569e1;
assign v855acb = EMPTY_p & v88ab6c | !EMPTY_p & v8a3239;
assign v8562d8 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8711d9;
assign v8a31b8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v856678;
assign BtoS_ACK1_n = !v85edf1;
assign v8550a0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855016;
assign v856bea = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v844f91;
assign v85579f = ENQ_p & v844fa9 | !ENQ_p & !v855d7f;
assign v86a9dc = RtoB_ACK0_p & v8563a6 | !RtoB_ACK0_p & v854ffa;
assign v8a3031 = jx0_p & v8a3194 | !jx0_p & v8a328d;
assign v860093 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v86aa63;
assign v856144 = EMPTY_p & v856723 | !EMPTY_p & v8563d8;
assign v8a2da1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v854d35;
assign v85621e = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & !v8a247a;
assign v855d2c = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v85e22c;
assign v8a333c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8a3334;
assign v8a3117 = EMPTY_p & v8558d2 | !EMPTY_p & v8a3062;
assign v856489 = jx2_p & v8a3222 | !jx2_p & v8a2cbd;
assign v8a3129 = StoB_REQ1_p & v855311 | !StoB_REQ1_p & v844f91;
assign v855e0d = jx1_p & v844f91 | !jx1_p & v8a329d;
assign v854eff = jx2_p & v8549bd | !jx2_p & !v85685d;
assign v8a311e = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v8a2f7a;
assign v855501 = jx2_p & v87119a | !jx2_p & v844f91;
assign v8a30b2 = StoB_REQ1_p & v8a30de | !StoB_REQ1_p & v844f91;
assign v8a336d = StoB_REQ1_p & v855e66 | !StoB_REQ1_p & v844f91;
assign v8a2fa9 = stateG7_1_p & v873756 | !stateG7_1_p & v844f91;
assign v844fbd = ENQ_p & v844f91 | !ENQ_p & !v844f91;
assign v8a29e3 = StoB_REQ1_p & v8551d0 | !StoB_REQ1_p & v844f91;
assign v856af3 = BtoS_ACK2_p & v844fa0 | !BtoS_ACK2_p & v856562;
assign v8a30c4 = DEQ_p & v8a3286 | !DEQ_p & v87734d;
assign v8560c6 = StoB_REQ1_p & v867273 | !StoB_REQ1_p & v85754a;
assign v8a3158 = jx0_p & v856e00 | !jx0_p & v8a31b3;
assign v855e40 = jx0_p & v854feb | !jx0_p & v8a3290;
assign v8a2fd5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v8a3187 = EMPTY_p & v844f91 | !EMPTY_p & v855af2;
assign v85685d = jx1_p & v8a3399 | !jx1_p & !v8a315a;
assign v855df9 = jx1_p & v8a2489 | !jx1_p & v896275;
assign v854f2f = ENQ_p & v8a3211 | !ENQ_p & v8a329f;
assign v855298 = jx2_p & v856835 | !jx2_p & v855254;
assign v8559ee = BtoS_ACK0_p & v856ab3 | !BtoS_ACK0_p & v85544e;
assign v856434 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85aae3;
assign v8562b9 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v8a31a7;
assign v86f89c = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8575b3;
assign v854ba4 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v873869;
assign v8a307c = ENQ_p & v856c57 | !ENQ_p & v8a3405;
assign v8a339d = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v877887;
assign v8a309d = stateG7_1_p & v8a30dd | !stateG7_1_p & v8a30e0;
assign v856c80 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v855c3e;
assign v8557be = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v888ecd;
assign v856871 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a313a;
assign v8a3393 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v8679b5 = BtoS_ACK1_p & v854b7c | !BtoS_ACK1_p & !v857619;
assign v8556cb = FULL_p & v85759c | !FULL_p & v855f60;
assign v854b14 = jx0_p & v856c72 | !jx0_p & v844f91;
assign SLC0_n = !v8961d4;
assign v8a3389 = StoB_REQ1_p & v85586d | !StoB_REQ1_p & v844f91;
assign v86aa49 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a316d;
assign jx1_n = !v866887;
assign v855fec = RtoB_ACK0_p & v855845 | !RtoB_ACK0_p & v856ab0;
assign v857a54 = StoB_REQ0_p & v8a31a7 | !StoB_REQ0_p & !v844f91;
assign v88ac3b = DEQ_p & v883c9a | !DEQ_p & v856c36;
assign v8a3086 = StoB_REQ3_p & v844f9f | !StoB_REQ3_p & v844f91;
assign v856bd6 = BtoS_ACK0_p & v87c725 | !BtoS_ACK0_p & v855ff1;
assign v8a283c = jx0_p & v856885 | !jx0_p & v844f91;
assign v8569e1 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v85581e;
assign v8a3405 = jx2_p & v856ad5 | !jx2_p & !v8a304d;
assign v873866 = RtoB_ACK1_p & v8a3293 | !RtoB_ACK1_p & v88ab9b;
assign v88abaa = stateG7_1_p & v8a2ef9 | !stateG7_1_p & v855ac2;
assign v85566d = DEQ_p & v856828 | !DEQ_p & v86dd6d;
assign v8a3289 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v85522d;
assign v8a300d = jx0_p & v8a312b | !jx0_p & !v857a21;
assign v8711ac = jx1_p & v856926 | !jx1_p & v854cc4;
assign v8a304e = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8576d5;
assign v85623b = FULL_p & v856432 | !FULL_p & v8a307b;
assign v8552b4 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v85555c;
assign v85a3a7 = BtoS_ACK1_p & v86c421 | !BtoS_ACK1_p & v896107;
assign v8a331e = jx0_p & v8a3355 | !jx0_p & v8a3249;
assign v8a3211 = jx2_p & v86f537 | !jx2_p & !v844f91;
assign v8a317f = jx1_p & v8961ac | !jx1_p & !v8a284d;
assign v856e10 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v8564c9;
assign v85555c = StoB_REQ3_p & v8a3315 | !StoB_REQ3_p & !v85523e;
assign v8a3235 = BtoS_ACK0_p & v844f9d | !BtoS_ACK0_p & v86a9cb;
assign v857651 = StoB_REQ0_p & v8550f3 | !StoB_REQ0_p & v8560bc;
assign v855894 = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v855600;
assign v856670 = BtoS_ACK0_p & v8711c0 | !BtoS_ACK0_p & v8a2d1f;
assign v8a33c6 = jx0_p & v855858 | !jx0_p & !v844f91;
assign v8a3178 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v856bc0;
assign v88abc1 = EMPTY_p & v857a8c | !EMPTY_p & v8557cd;
assign v88ab43 = ENQ_p & v87c729 | !ENQ_p & v857418;
assign v8a3244 = jx2_p & v8a33ae | !jx2_p & v856e3f;
assign v857521 = StoB_REQ2_p & v856e2b | !StoB_REQ2_p & v8a243e;
assign v8550fb = BtoS_ACK0_p & v8562d8 | !BtoS_ACK0_p & v8a2da1;
assign v8554bf = BtoS_ACK1_p & v8711c0 | !BtoS_ACK1_p & v8617be;
assign v87119a = jx1_p & v844f91 | !jx1_p & !v855cb6;
assign v8a314b = StoB_REQ2_p & v8a29a5 | !StoB_REQ2_p & v8a3354;
assign v857547 = jx0_p & v856670 | !jx0_p & v8a321d;
assign v85741f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v855f5b;
assign v8a31fe = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v855042;
assign v8a2c62 = stateG7_1_p & v85500c | !stateG7_1_p & v8a3131;
assign v85679c = BtoR_REQ1_p & v8a31fd | !BtoR_REQ1_p & v86d760;
assign v8560ea = BtoS_ACK4_p & v844f9d | !BtoS_ACK4_p & !v844f91;
assign v854204 = DEQ_p & v8a31af | !DEQ_p & v8a30be;
assign v8558f4 = StoB_REQ0_p & v8565b9 | !StoB_REQ0_p & v844f91;
assign v86b201 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a3268;
assign v85614f = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v854b5f;
assign v855047 = EMPTY_p & v855ead | !EMPTY_p & v8a3304;
assign v896162 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855533;
assign v855033 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a312e;
assign v8a30e9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v85614f;
assign v855631 = jx0_p & v8574ee | !jx0_p & v844f9d;
assign v8a2b19 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v854c82;
assign v8558cb = EMPTY_p & v8a32c6 | !EMPTY_p & v8a2486;
assign v8685f8 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & !v8a336c;
assign v8a30b0 = jx1_p & v856786 | !jx1_p & v8a3245;
assign v855fb0 = ENQ_p & v8a317d | !ENQ_p & v844f91;
assign v857689 = DEQ_p & v8a338e | !DEQ_p & v8556cb;
assign v854d01 = jx1_p & v844f91 | !jx1_p & v85747f;
assign v855c3a = StoB_REQ0_p & v8a2b16 | !StoB_REQ0_p & v857a0c;
assign v85ecec = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v8a30b3;
assign v87116e = stateG7_1_p & v8a3228 | !stateG7_1_p & v855ea7;
assign v854ed7 = ENQ_p & v8a313f | !ENQ_p & v856847;
assign v8a247a = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v8a31bd;
assign v8a2c6b = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v844f9d;
assign v8a3040 = DEQ_p & v85786a | !DEQ_p & v86dd6d;
assign v8a3282 = StoB_REQ0_p & v8550f3 | !StoB_REQ0_p & v856863;
assign v8a2e00 = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & v88b745;
assign v854fc7 = ENQ_p & v87bbfb | !ENQ_p & v876345;
assign v8a30a5 = jx1_p & v855a2a | !jx1_p & v844fa9;
assign v8a28a9 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v8a30dc;
assign v8a3176 = jx0_p & v8a3260 | !jx0_p & !v8617fe;
assign v85743c = DEQ_p & v8a3058 | !DEQ_p & !v854fc1;
assign v8a3147 = StoB_REQ2_p & v8a283f | !StoB_REQ2_p & v844f91;
assign v8532c4 = StoB_REQ3_p & v854ee4 | !StoB_REQ3_p & v844f91;
assign v8574ee = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v8a2893;
assign jx0_n = !v8711df;
assign v856cd1 = stateG12_p & v85613d | !stateG12_p & !v844f91;
assign v8a29ad = BtoS_ACK0_p & v844f9f | !BtoS_ACK0_p & v854b33;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v855eb2 = StoB_REQ2_p & v844f9d | !StoB_REQ2_p & v844f91;
assign v868cba = BtoS_ACK0_p & v855fdf | !BtoS_ACK0_p & !v8a30b4;
assign v8a33df = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v855e1c;
assign v855833 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v855ef6;
assign v844fa1 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v88a469 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8558f4;
assign v856062 = StoB_REQ2_p & v856acb | !StoB_REQ2_p & v8a31c1;
assign v857a21 = BtoS_ACK0_p & v854a11 | !BtoS_ACK0_p & v8a31e2;
assign v856bdb = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v855531;
assign v856705 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v861796;
assign v854b1e = StoB_REQ2_p & v844f9f | !StoB_REQ2_p & v876d51;
assign v88abed = BtoS_ACK0_p & v8711cf | !BtoS_ACK0_p & v8a336a;
assign v86b41a = jx2_p & v8a31f4 | !jx2_p & v85617a;
assign v8551ba = DEQ_p & v8a338e | !DEQ_p & v8a3049;
assign v8565b9 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v8555ef;
assign v855c5f = StoB_REQ1_p & v85699f | !StoB_REQ1_p & v856e5f;
assign v857414 = EMPTY_p & v855d44 | !EMPTY_p & v8962f6;
assign v8a2b13 = DEQ_p & v8554e5 | !DEQ_p & v85623b;
assign v88ab87 = BtoS_ACK1_p & v844fa0 | !BtoS_ACK1_p & v8a3132;
assign v8a3166 = StoB_REQ2_p & v8a331b | !StoB_REQ2_p & v854d33;
assign v8a3303 = StoB_REQ3_p & v854f52 | !StoB_REQ3_p & v857731;
assign v88a46b = StoB_REQ2_p & v855033 | !StoB_REQ2_p & v8a339d;
assign v8a2bf7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v854e7c;
assign v85749f = BtoR_REQ1_p & v8961cb | !BtoR_REQ1_p & v8960ee;
assign v8a3364 = EMPTY_p & v856723 | !EMPTY_p & v8551ba;
assign v873899 = StoB_REQ3_p & v854f52 | !StoB_REQ3_p & v85523e;
assign v854ee4 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844f9f;
assign v856df1 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v8a30ac;
assign v85663b = BtoS_ACK0_p & v8711c0 | !BtoS_ACK0_p & v8a3229;
assign v855cb6 = jx0_p & v8a312b | !jx0_p & !v844f91;
assign v86f537 = jx1_p & v844f91 | !jx1_p & !v844f91;
assign v8a33cd = BtoS_ACK0_p & v856c06 | !BtoS_ACK0_p & v856e26;
assign v857932 = BtoS_ACK0_p & v8a2972 | !BtoS_ACK0_p & v861d68;
assign v88ab71 = StoB_REQ0_p & v8774cb | !StoB_REQ0_p & v855a89;
assign v8a2f81 = ENQ_p & v856c57 | !ENQ_p & v8574f8;
assign v854a71 = StoB_REQ3_p & v854bf7 | !StoB_REQ3_p & v857731;
assign v8566ad = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a3358;
assign v8a2935 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v8a308c;
assign v8558cf = BtoS_ACK0_p & v855c79 | !BtoS_ACK0_p & v85677d;
assign v8a3220 = StoB_REQ0_p & v8553e6 | !StoB_REQ0_p & v8738ae;
assign v8a31bd = BtoS_ACK4_p & v844f91 | !BtoS_ACK4_p & v844f9d;
assign v8a33ce = StoB_REQ2_p & v8a3082 | !StoB_REQ2_p & v8a2d78;
assign v854a65 = StoB_REQ0_p & v8774cb | !StoB_REQ0_p & v855d54;
assign v8a2f21 = BtoS_ACK5_p & v844f91 | !BtoS_ACK5_p & v844f9f;
assign v855aec = StoB_REQ0_p & v8a30b1 | !StoB_REQ0_p & v844f91;
assign v8a32df = BtoS_ACK0_p & v856883 | !BtoS_ACK0_p & v8a31d2;
assign v856db6 = BtoR_REQ1_p & v8a2e76 | !BtoR_REQ1_p & v855a4d;
assign v867269 = jx2_p & v8a2e8b | !jx2_p & v856b69;
assign v85edc7 = StoB_REQ3_p & v86aa63 | !StoB_REQ3_p & v844fb1;
assign v87d011 = BtoS_ACK1_p & v854b1e | !BtoS_ACK1_p & v8a33c7;
assign v8a32c0 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a3207;
assign v8a2bb0 = jx2_p & v85ed1a | !jx2_p & !v8a30ce;
assign v8a31f3 = StoB_REQ0_p & v855600 | !StoB_REQ0_p & v856bdb;
assign v85a4b2 = jx0_p & v856966 | !jx0_p & v844f91;
assign v8a2f08 = FULL_p & v8541c7 | !FULL_p & v8a3048;
assign v8557b8 = BtoS_ACK0_p & v8a32f4 | !BtoS_ACK0_p & v8a3099;
assign v8a3091 = jx1_p & v8a2fd5 | !jx1_p & v855870;
assign v8a3309 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v8a31d8;
assign v8a29d7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v8a31ca;
assign v854f98 = stateG7_1_p & v855b1d | !stateG7_1_p & v857775;
assign v8a2d5b = jx0_p & v854c5b | !jx0_p & !v8a24a6;
assign v8a31e6 = EMPTY_p & v855d44 | !EMPTY_p & v855fb5;
assign v856885 = BtoS_ACK0_p & v855c79 | !BtoS_ACK0_p & v854a65;
assign v856102 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v8553de;
assign v8a32eb = StoB_REQ1_p & v8a29d7 | !StoB_REQ1_p & v8a333c;
assign v854c99 = jx1_p & v856786 | !jx1_p & v8a3206;
assign v8a308f = ENQ_p & v844f91 | !ENQ_p & v8a3154;
assign v8559bc = EMPTY_p & v856063 | !EMPTY_p & v8a32fb;
assign v8a3391 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a3393;
assign v856e02 = stateG7_1_p & v883cae | !stateG7_1_p & v861800;
assign v89caa5 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v856062;
assign v8a309b = jx2_p & v85e7e0 | !jx2_p & v8711ac;
assign v8a31c1 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v855790;
assign v855314 = jx2_p & v87c300 | !jx2_p & !v8a30e2;
assign v8a3380 = jx1_p & v85606a | !jx1_p & v8a325f;
assign v8711df = BtoR_REQ0_p & v8a3288 | !BtoR_REQ0_p & v85749f;
assign v8a32b8 = jx2_p & v856575 | !jx2_p & !v8a31ea;
assign v8a3321 = BtoR_REQ1_p & v8a328e | !BtoR_REQ1_p & v856256;
assign v8a32d7 = EMPTY_p & v8a2f81 | !EMPTY_p & !v8a31bc;
assign v855114 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v8a3303;
assign v8a322d = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v85532e;
assign v8960fd = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a315b;
assign SLC1_n = !v88a46f;
assign v8563a6 = EMPTY_p & v87c707 | !EMPTY_p & v855cfe;
assign v856926 = jx0_p & v8a3258 | !jx0_p & v8960fd;
assign v85683b = ENQ_p & v855298 | !ENQ_p & v85508c;
assign v8576d5 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v8a30b2;
assign v88abca = jx1_p & v8573f3 | !jx1_p & v85741f;
assign v8711cf = StoB_REQ1_p & v844f9d | !StoB_REQ1_p & v85ed6f;
assign v855d6a = BtoS_ACK0_p & v857969 | !BtoS_ACK0_p & v8a30c5;
assign v85523e = StoB_REQ4_p & v844f9f | !StoB_REQ4_p & v844f91;
assign v86aa4a = EMPTY_p & v8a2984 | !EMPTY_p & v8a3304;
assign v856a09 = BtoS_ACK1_p & v856639 | !BtoS_ACK1_p & v8a3395;
assign v8a3189 = jx1_p & v856b69 | !jx1_p & v8a2d89;
assign v8579f3 = BtoS_ACK0_p & v8a336d | !BtoS_ACK0_p & v8a3285;
assign v87116b = BtoS_ACK2_p & v844f9d | !BtoS_ACK2_p & v854a11;
assign v8a317d = jx2_p & v855ddf | !jx2_p & v856553;
assign v8566b6 = jx2_p & v844f91 | !jx2_p & v8a0e3c;
assign v8a2485 = StoB_REQ2_p & v8a331b | !StoB_REQ2_p & v8a33b2;
assign v8a3052 = jx1_p & v8a3151 | !jx1_p & v8a3176;
assign v8a30ac = StoB_REQ2_p & v8a283f | !StoB_REQ2_p & v8552f8;
assign v854a17 = BtoS_ACK1_p & v8a337f | !BtoS_ACK1_p & v854a89;
assign v8a32d0 = EMPTY_p & v876d41 | !EMPTY_p & v855a61;
assign v8a28af = DEQ_p & v856901 | !DEQ_p & v856063;
assign v85532e = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & v844f9d;
assign v85634e = BtoS_ACK1_p & v8a3032 | !BtoS_ACK1_p & v8a32eb;
assign v856648 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v85540d;
assign v865746 = ENQ_p & v86178d | !ENQ_p & v8a2ee2;
assign v8a304c = jx2_p & v854d3e | !jx2_p & v85606a;
assign v85786a = ENQ_p & v8a302e | !ENQ_p & !v855d7f;
assign v856130 = stateG7_1_p & v8a30ab | !stateG7_1_p & v8550c7;
assign v8a31c7 = jx2_p & v8a3052 | !jx2_p & v8555a0;
assign v8556ec = DEQ_p & v8a3058 | !DEQ_p & !v8a2c65;
assign v8a3095 = jx2_p & v8a33ac | !jx2_p & !v8a304d;
assign v87c76f = BtoR_REQ0_p & v857b8b | !BtoR_REQ0_p & v85e12c;
assign v85644e = StoB_REQ1_p & v854b5f | !StoB_REQ1_p & v856352;
assign v8a31ed = BtoS_ACK3_p & v844f9d | !BtoS_ACK3_p & v8a31bd;
assign v8a33b0 = jx2_p & v87119a | !jx2_p & !v855df9;
assign v8a3253 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v85586a;
assign v8a2fe8 = StoB_REQ0_p & v8774cb | !StoB_REQ0_p & v854eb2;
assign v8a338c = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855cd0;
assign v856374 = jx0_p & v856781 | !jx0_p & v8a2fba;
assign v8a3229 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8567b5;
assign v85d977 = ENQ_p & v855254 | !ENQ_p & v8a32ce;
assign v8a0e0a = StoB_REQ1_p & v8630d3 | !StoB_REQ1_p & v8a3115;
assign v856835 = jx1_p & v855254 | !jx1_p & v85796e;
assign v855fac = DEQ_p & v8a30a6 | !DEQ_p & v85651f;
assign v857a31 = StoB_REQ1_p & v8a2972 | !StoB_REQ1_p & v854b1e;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v854a06 = jx1_p & v856624 | !jx1_p & !v8a3372;
assign v86938f = StoB_REQ0_p & v8961a8 | !StoB_REQ0_p & v857aed;
assign v855078 = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v856636;
assign v896248 = StoB_REQ0_p & v85eb80 | !StoB_REQ0_p & v855c86;
assign v8a3049 = ENQ_p & v8574eb | !ENQ_p & v85660e;
assign v8a327e = DEQ_p & v883c9a | !DEQ_p & v85797a;
assign v8551d0 = BtoS_ACK2_p & v844f9b | !BtoS_ACK2_p & v8a3350;
assign v854be5 = jx0_p & v8a30e7 | !jx0_p & !v85698e;
assign v857534 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a32c4;
assign v8a329c = ENQ_p & v856553 | !ENQ_p & v844f91;
assign v855196 = jx1_p & v8a3313 | !jx1_p & v854be5;
assign v8556a7 = EMPTY_p & v854fcb | !EMPTY_p & !v854fc7;
assign v8617fe = BtoS_ACK0_p & v854a11 | !BtoS_ACK0_p & v854ffe;
assign v854c82 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v871051;
assign v856992 = DEQ_p & v8a3058 | !DEQ_p & v844f91;
assign v854cbb = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3225;
assign v855d7f = jx2_p & v8a310a | !jx2_p & v8711ac;
assign v8a3033 = StoB_REQ1_p & v8a3314 | !StoB_REQ1_p & v86aa4d;
assign v8a332e = BtoS_ACK1_p & v88ab81 | !BtoS_ACK1_p & v8a29d7;
assign v854ae3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a32a4;
assign v8617be = BtoS_ACK2_p & v8a3086 | !BtoS_ACK2_p & v88a46b;
assign v8a330a = ENQ_p & v8a324a | !ENQ_p & v8a3030;
assign v855d7a = jx0_p & v85528e | !jx0_p & !v8562b9;
assign v855b5d = EMPTY_p & v854d31 | !EMPTY_p & v855cc1;
assign v8a3206 = jx0_p & v855bdb | !jx0_p & v856431;
assign v856b2a = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v85754a;
assign v8a3107 = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v855db1;
assign v8a2f6b = BtoS_ACK1_p & v8a337f | !BtoS_ACK1_p & v857af8;
assign v8a2cab = BtoS_ACK3_p & v855b05 | !BtoS_ACK3_p & v857692;
assign v85797a = FULL_p & v856432 | !FULL_p & v85651f;
assign v8558fe = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v855ef6;
assign v854c39 = stateG7_1_p & v86aa3d | !stateG7_1_p & v89614f;
assign v861784 = BtoS_ACK2_p & v844f9f | !BtoS_ACK2_p & v854c5c;
assign v8a3314 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v8a3082;
assign v8a3088 = FULL_p & v844f91 | !FULL_p & v85640f;
assign v85577c = BtoS_ACK0_p & v856c06 | !BtoS_ACK0_p & v8a2b42;
assign v8573f3 = stateG12_p & v85741f | !stateG12_p & v844f91;
assign v856e7f = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v872af1;
assign v855ebc = jx1_p & v85698e | !jx1_p & !v8a320a;
assign v8a3208 = StoB_REQ0_p & v8573cd | !StoB_REQ0_p & v855e0e;
assign v855397 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3178;
assign v8a307a = jx2_p & v8a297d | !jx2_p & !v844f91;
assign v844fbf = DEQ_p & v844f91 | !DEQ_p & !v844f91;
assign v8a3350 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v855ef6;
assign v854c76 = BtoS_ACK4_p & v869886 | !BtoS_ACK4_p & v8a2f21;
assign v8a3330 = BtoS_ACK1_p & v855311 | !BtoS_ACK1_p & !v873869;
assign v8a324c = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v857534;
assign v857421 = StoB_REQ1_p & v86f89c | !StoB_REQ1_p & v8a3023;
assign v8a2c6e = ENQ_p & v844fa9 | !ENQ_p & !v85528a;
assign v8a30d1 = jx2_p & v856b4c | !jx2_p & !v8703da;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v8a3267 = RtoB_ACK1_p & v857572 | !RtoB_ACK1_p & v8a3397;
assign v8a32a4 = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v8a3096;
assign v856c72 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v85618d;
assign v855283 = DEQ_p & v8a31af | !DEQ_p & v855f60;
assign v855708 = StoB_REQ0_p & v844f9d | !StoB_REQ0_p & v8a2ff0;
assign v8a33c4 = jx2_p & v854d3e | !jx2_p & v844f91;
assign v8a3246 = StoB_REQ1_p & v8562d8 | !StoB_REQ1_p & v844f91;
assign v857a0c = BtoS_ACK1_p & v85ed6f | !BtoS_ACK1_p & v8560c6;
assign v8a3258 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v855edf;
assign v883754 = EMPTY_p & v854ed7 | !EMPTY_p & v8a31e5;
assign v85a137 = ENQ_p & v8a324a | !ENQ_p & v855314;
assign v855414 = EMPTY_p & v856b58 | !EMPTY_p & v8961a7;
assign v85594d = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8579fd;
assign v856b26 = jx2_p & v86eb76 | !jx2_p & v85413e;
assign v8553cf = BtoS_ACK1_p & v844f9d | !BtoS_ACK1_p & v8558d9;
assign v855147 = StoB_REQ0_p & v8774cb | !StoB_REQ0_p & v856313;
assign v8a31b1 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a3307;
assign v88abdb = StoB_REQ1_p & v854b5f | !StoB_REQ1_p & v8a3135;
assign v856497 = jx1_p & v844f91 | !jx1_p & v855739;
assign v873280 = jx1_p & v844fc1 | !jx1_p & v844f91;
assign v855e0c = ENQ_p & v856b26 | !ENQ_p & v8a2b44;
assign v856075 = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v8568b1;
assign v8a30ec = DEQ_p & v8a3058 | !DEQ_p & !v86cbc9;
assign v8552ea = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v854e78;
assign v8a30cf = ENQ_p & v85610f | !ENQ_p & v858bbc;
assign v8567c7 = StoB_REQ3_p & v856d89 | !StoB_REQ3_p & v844f91;
assign v8a3144 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v86f804;
assign v85793b = jx1_p & v8a3156 | !jx1_p & !v85646a;
assign v8a3115 = BtoS_ACK2_p & v8a3036 | !BtoS_ACK2_p & v8a2e9b;
assign v8a30e0 = EMPTY_p & v8a3221 | !EMPTY_p & v855283;
assign v855fb5 = DEQ_p & v896289 | !DEQ_p & v8a329c;
assign v8579fd = BtoS_ACK1_p & v855eb2 | !BtoS_ACK1_p & v8a31ac;
assign v856aa1 = jx2_p & v8541c3 | !jx2_p & v8a326b;
assign v855b05 = StoB_REQ4_p & v844f91 | !StoB_REQ4_p & v844fa0;
assign v85509f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8a320d;
assign v856e34 = StoB_REQ1_p & v855a7a | !StoB_REQ1_p & v8a30fd;
assign v8a3222 = jx1_p & v844fc1 | !jx1_p & !v8a33db;
assign v8a318a = BtoS_ACK1_p & v856639 | !BtoS_ACK1_p & v8a0e0a;
assign v855653 = jx2_p & v8a2e72 | !jx2_p & v855254;
assign v8711bb = EMPTY_p & v844f91 | !EMPTY_p & v8a3236;
assign v854fff = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a2d93;
assign v8a2898 = EMPTY_p & v857649 | !EMPTY_p & v88ac3b;
assign v8a313a = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v8a3354;
assign v85499f = jx0_p & v85413d | !jx0_p & v8a0de9;
assign v888edb = BtoR_REQ0_p & v8549ca | !BtoR_REQ0_p & v856c11;
assign v88a44b = BtoS_ACK2_p & v876d51 | !BtoS_ACK2_p & v8a31cd;
assign v857b8b = RtoB_ACK0_p & v857a7a | !RtoB_ACK0_p & v856130;
assign v8a3345 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8a3305;
assign v85751a = BtoS_ACK1_p & v844f9f | !BtoS_ACK1_p & v87d020;
assign v856b58 = ENQ_p & v855254 | !ENQ_p & v855709;
assign v8a3043 = jx0_p & v856aac | !jx0_p & v844f91;
assign v85681c = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v8a3186;
assign v883730 = BtoS_ACK3_p & v844f9f | !BtoS_ACK3_p & !v8a336c;
assign v8a32d8 = stateG7_1_p & v8a3171 | !stateG7_1_p & v88abc1;
assign v8a2d0e = ENQ_p & v844f91 | !ENQ_p & v855501;
assign ENQ_n = (stateG7_1_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((StoB_REQ0_n))) | (!jx1_n & ((jx0_n) | (!jx0_n & ((StoB_REQ0_n))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))))))))))) | (!stateG7_0_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((jx2_n) | (!jx2_n & ((jx1_n) | (!jx1_n & ((jx0_n))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((StoB_REQ0_n))) | (!jx1_n & ((jx0_n) | (!jx0_n & ((StoB_REQ0_n))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))) | (!jx0_n & ((BtoS_ACK1_n) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!DEQ_n & ((stateG12_n & ((!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n))))))))))))))))) | (!stateG12_n & ((!FULL_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((StoB_REQ2_n))) | (!BtoS_ACK2_n & ((SLC1_n & ((!SLC2_n & ((SLC0_n))))) | (!SLC1_n & ((SLC2_n) | (!SLC2_n & ((SLC0_n)))))))))))))))))))))))))));
assign SLC2_n = (stateG7_1_n & ((stateG7_0_n & ((BtoR_REQ0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!jx1_n & ((!jx0_n & ((!StoB_REQ0_n & ((SLC1_n))))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!jx1_n & ((!jx0_n & ((!StoB_REQ0_n & ((SLC1_n))))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))))) | (!stateG7_0_n & ((BtoR_REQ0_n & ((RtoB_ACK0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK0_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!jx1_n & ((!jx0_n & ((!StoB_REQ0_n & ((SLC1_n))))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((RtoB_ACK1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))) | (!RtoB_ACK1_n & ((EMPTY_n & ((jx2_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!jx2_n & ((!BtoS_ACK0_n & ((jx1_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))) | (!jx1_n & ((jx0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))))))))))) | (!stateG7_1_n & ((BtoR_REQ0_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!BtoR_REQ0_n & ((RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((!SLC1_n))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!StoB_REQ1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))) | (!StoB_REQ2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((StoB_REQ3_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))) | (!StoB_REQ3_n & ((SLC0_n))))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))))))))) | (!RtoB_ACK0_n & ((BtoR_REQ1_n & ((EMPTY_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))))) | (!BtoR_REQ1_n & ((EMPTY_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((!BtoS_ACK3_n))) | (!SLC1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((jx1_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!jx1_n & ((!jx0_n & ((!StoB_REQ0_n & ((SLC1_n))))))))) | (!BtoS_ACK0_n & ((jx1_n & ((jx0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))) | (!jx0_n & ((!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!EMPTY_n & ((DEQ_n & ((stateG12_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))) | (!stateG12_n & ((SLC1_n))))) | (!DEQ_n & ((stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((!BtoS_ACK3_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))) | (!jx1_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))) | (!jx2_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n))))))))))))))))))))) | (!stateG12_n & ((FULL_n & ((SLC1_n))) | (!FULL_n & ((BtoS_ACK0_n & ((!StoB_REQ0_n & ((SLC1_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((!StoB_REQ1_n & ((SLC1_n))))) | (!BtoS_ACK1_n & ((BtoS_ACK2_n & ((!StoB_REQ2_n & ((SLC1_n))))) | (!BtoS_ACK2_n & ((SLC1_n & ((StoB_REQ3_n & ((!BtoS_ACK3_n))) | (!StoB_REQ3_n))) | (!SLC1_n & ((BtoS_ACK3_n & ((SLC0_n))) | (!BtoS_ACK3_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ4_n & ((BtoS_ACK4_n)))))))))))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  StoB_REQ4_p = 0;
  StoB_REQ5_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoS_ACK4_p = 0;
  BtoS_ACK5_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  SLC2_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  StoB_REQ4_p = StoB_REQ4_n;
  StoB_REQ5_p = StoB_REQ5_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoS_ACK4_p = BtoS_ACK4_n;
  BtoS_ACK5_p = BtoS_ACK5_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  SLC2_p = SLC2_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
