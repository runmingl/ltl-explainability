module main(clock, StoB_REQ0_n, StoB_REQ1_n, StoB_REQ2_n, StoB_REQ3_n, RtoB_ACK0_n, RtoB_ACK1_n, FULL_n, EMPTY_n, BtoS_ACK0_n, BtoS_ACK1_n, BtoS_ACK2_n, BtoS_ACK3_n, BtoR_REQ0_n, BtoR_REQ1_n, stateG7_0_n, stateG7_1_n, ENQ_n, DEQ_n, stateG12_n, SLC0_n, SLC1_n, jx0_n, jx1_n, jx2_n);
  input clock;
  wire zero_value = 0;
  wire one_value = 1;
  wire v844f91;
  wire v844f99;
  wire v873071;
  wire v87eca7;
  wire v872dd8;
  wire v87eef6;
  wire v8733ec;
  wire v85b574;
  wire v87eda4;
  wire v8582c0;
  wire v868b92;
  wire v87ecd5;
  wire v873774;
  wire v87377f;
  wire v844f9b;
  wire v859947;
  wire v872ee2;
  wire v87ede2;
  wire v872da9;
  wire v87edcc;
  wire v87eccc;
  wire v844fad;
  wire v844f9f;
  wire v87283c;
  wire v872d64;
  wire v87edc4;
  wire v872d99;
  wire v872878;
  wire v8757d4;
  wire v87edb2;
  wire v87e848;
  wire v87372e;
  wire v876322;
  wire v872835;
  wire v87ed06;
  wire v8750bd;
  wire v874051;
  wire v87ec1b;
  wire v87ecda;
  wire v87e8e1;
  wire v87305a;
  wire v872fa1;
  wire v872e0f;
  wire v873172;
  wire v8737e3;
  wire v87eee0;
  wire v858b3f;
  wire v87edc6;
  wire v873078;
  wire v87ec49;
  wire v87ecea;
  wire v872f13;
  wire v872ee9;
  wire v868baa;
  wire v873784;
  wire v872df4;
  wire v87ebe9;
  wire v862858;
  wire v844fb3;
  wire v87edcb;
  wire v87ed9f;
  wire v87ec2d;
  wire v85409b;
  wire v852e67;
  wire v8732d3;
  wire v87ec9f;
  wire v872c60;
  wire v87ed62;
  wire v872c81;
  wire v872e9a;
  wire v872b5c;
  wire v87ecd7;
  wire v87ec12;
  wire v87ed1e;
  wire v87ed79;
  wire v87ebee;
  wire v87378d;
  wire v87ee84;
  wire v872949;
  wire v872fbc;
  wire v87ed51;
  wire v8733af;
  wire v858bae;
  wire v87ee0f;
  wire v87ec72;
  wire v87ec51;
  wire v873370;
  wire v855cab;
  wire v87efc9;
  wire v87efc2;
  wire v874df5;
  wire v872e81;
  wire v876314;
  wire v85abe7;
  wire v872d4f;
  wire v85271e;
  wire v875111;
  wire v8733e9;
  wire v852d87;
  wire v872fa7;
  wire v8732c4;
  wire v873327;
  wire v87ec05;
  wire v876307;
  wire v874bf2;
  wire v8752b0;
  wire v872d6b;
  wire v8757d7;
  wire v872fb8;
  wire v87eeaa;
  wire v87338a;
  wire v87ebe4;
  wire v8598e6;
  wire v87ec5a;
  wire v87ec96;
  wire v8731d4;
  wire v87eceb;
  wire v87efce;
  wire v85448e;
  wire v873079;
  wire v874c38;
  wire v872877;
  wire v87ed8f;
  wire v87ec28;
  wire v872de4;
  wire v87eda9;
  wire v87ed80;
  wire v87ecc6;
  wire v872f69;
  wire v8745a9;
  wire v87edd7;
  wire v872dbf;
  wire v8567f5;
  wire v8728e2;
  wire v87ed27;
  wire v879395;
  wire v85b5e0;
  wire v844faf;
  wire v873197;
  wire v872f4e;
  wire v86e02d;
  wire v87ec2c;
  wire v8745a5;
  wire v854111;
  wire v87307b;
  wire v87ed3d;
  wire v87ecef;
  wire v87ecd2;
  wire v872db6;
  wire v87ed0b;
  wire v87ec0b;
  wire v87622d;
  wire v87ed75;
  wire v872c19;
  wire v856719;
  wire v873307;
  wire v87eddd;
  wire v8728a3;
  wire v87ecbf;
  wire v8727f7;
  wire v872ec6;
  wire v876238;
  wire v853052;
  wire v8757c5;
  wire v86283e;
  wire v872f60;
  wire v87e8f1;
  wire v872f1a;
  wire v8589e8;
  wire v87ec7a;
  wire v87ebfe;
  wire v872ec1;
  wire v87e85d;
  wire v872fa5;
  wire v8728d6;
  wire v87ed5b;
  wire v87ec5e;
  wire v852d6f;
  wire v87ec1a;
  wire v876245;
  wire v87379c;
  wire v872cd6;
  wire v87ec6b;
  wire v87ed7b;
  wire v855c35;
  wire v8588f4;
  wire v87ecd1;
  wire v87ed83;
  wire v87ed2f;
  wire v87ed84;
  wire v87e8f3;
  wire v87ed3f;
  wire v87ec0a;
  wire v872ec9;
  wire v872fee;
  wire v872c17;
  wire v87422b;
  wire v87eccf;
  wire v852626;
  wire v87ebf4;
  wire v87ec14;
  wire v872e92;
  wire v8757d2;
  wire v87ec95;
  wire v852227;
  wire v868b30;
  wire v85a741;
  wire v85a712;
  wire v853eb8;
  wire v87ec42;
  wire v868af3;
  wire v86284b;
  wire v87edb3;
  wire v8728c0;
  wire v8686b4;
  wire v872e99;
  wire v872d67;
  wire v85a0a4;
  wire v8752ab;
  wire v87ee02;
  wire v87ec19;
  wire v873077;
  wire v87ed47;
  wire v8730b0;
  wire v868b71;
  wire v872e80;
  wire v87623a;
  wire v852eb2;
  wire v87ed92;
  wire v87ef77;
  wire v873048;
  wire v872c93;
  wire v852d93;
  wire v872e09;
  wire v856f49;
  wire v868b8b;
  wire v87ec4a;
  wire v87ef9c;
  wire v857ea2;
  wire v872ed3;
  wire v87ed76;
  wire v87ec25;
  wire v874242;
  wire v872e6f;
  wire v8731c8;
  wire v87ecbd;
  wire v87ee8b;
  wire v872d7f;
  wire v87ed9d;
  wire v872f17;
  wire v87e8be;
  wire v87e82a;
  wire v87eda6;
  wire v87ed45;
  wire v87ecdb;
  wire v844f9d;
  wire v87ec41;
  wire v872f67;
  wire v8737c6;
  wire v872927;
  wire v87ef83;
  wire v87e855;
  wire v87e8df;
  wire v8728cb;
  wire v87eccb;
  wire v87ed13;
  wire v87287b;
  wire v87ec15;
  wire v872eb0;
  wire v872fe0;
  wire v8731b9;
  wire v872f47;
  wire v87302a;
  wire v8757c6;
  wire v873723;
  wire v872e8b;
  wire v87ed1c;
  wire v872819;
  wire v859541;
  wire v868ba1;
  wire v855989;
  wire v87322c;
  wire v87ec23;
  wire v87372a;
  wire v872f5d;
  wire v87e8d0;
  wire v85a673;
  wire v8733de;
  wire v87eca1;
  wire v87ec89;
  wire v858f67;
  wire v87ec98;
  wire v87ec1c;
  wire v87ef0a;
  wire v87ecfa;
  wire v8564be;
  wire v8737e4;
  wire v873333;
  wire v87ebf1;
  wire v858d4f;
  wire v873726;
  wire v868b3d;
  wire v87ed97;
  wire v87500a;
  wire v87e85b;
  wire v873177;
  wire v87291f;
  wire v868b4a;
  wire v87ebf5;
  wire v872f82;
  wire v872e7f;
  wire v85ab45;
  wire v872975;
  wire v87ec6d;
  wire v87ec53;
  wire v858bc4;
  wire v856718;
  wire v87323e;
  wire v87edd0;
  wire v87eec0;
  wire v87ed9e;
  wire v872dff;
  wire v872c51;
  wire v87ed48;
  wire v8730c6;
  wire v85b091;
  wire v87eca2;
  wire v8737ab;
  wire v87ec48;
  wire v85724c;
  wire v872bf1;
  wire v8730c8;
  wire v868ae0;
  wire v8572b7;
  wire v8594bd;
  wire v852226;
  wire v857f15;
  wire v85260c;
  wire v87332b;
  wire v87ec40;
  wire v8731a1;
  wire v868b9a;
  wire v87edf9;
  wire v8732f0;
  wire v872ecb;
  wire v872890;
  wire v87ee9d;
  wire v8731f8;
  wire v859412;
  wire v8733c1;
  wire v872e7a;
  wire v87ec06;
  wire v87ed10;
  wire v87370d;
  wire v873759;
  wire v872eae;
  wire v872e78;
  wire v868b6d;
  wire v87ecc3;
  wire v87ebef;
  wire v8757ca;
  wire v87318f;
  wire v8793a7;
  wire v873074;
  wire v872f4c;
  wire v872e22;
  wire v87ee95;
  wire v87ebe3;
  wire v8730f3;
  wire v872d03;
  wire v87ecb5;
  wire v87efcf;
  wire v872dca;
  wire v868b3a;
  wire v852d67;
  wire v87289c;
  wire v873392;
  wire v87edd5;
  wire v87332f;
  wire v87ecfd;
  wire v87ec11;
  wire v87ed96;
  wire v868adc;
  wire v87ecb6;
  wire v8525dc;
  wire v87ed23;
  wire v872e8e;
  wire v868bef;
  wire v844fb9;
  wire v87eee6;
  wire v879392;
  wire v87ec99;
  wire v872d56;
  wire v8737c4;
  wire v87330a;
  wire v844fab;
  wire v8750ad;
  wire v873799;
  wire v873293;
  wire v8733da;
  wire v868b29;
  wire v8736f4;
  wire v87ed3e;
  wire v874c37;
  wire v87ed01;
  wire v87ecbb;
  wire v872837;
  wire v8730eb;
  wire v85b2d3;
  wire v85adeb;
  wire v873741;
  wire v8731fb;
  wire v87ec32;
  wire v87ed61;
  wire v87ed04;
  wire v872936;
  wire v8731b2;
  wire v87ed36;
  wire v87ecde;
  wire v872b76;
  wire v868aba;
  wire v872f79;
  wire v868bde;
  wire v873176;
  wire v872ff7;
  wire v8538fd;
  wire v87bbdd;
  wire v87ec65;
  wire v87291a;
  wire v87ed70;
  wire v87ecb1;
  wire v87286f;
  wire v87ed3b;
  wire v87ed7a;
  wire v87ed6b;
  wire v87ec56;
  wire v8736f8;
  wire v873250;
  wire v87efcc;
  wire v87ec01;
  wire v872d35;
  wire v873375;
  wire v8728da;
  wire v872916;
  wire v857beb;
  wire v87ec71;
  wire v8732c2;
  wire v873779;
  wire v87ec8e;
  wire v87ebf6;
  wire v874064;
  wire v873379;
  wire v87e86b;
  wire v868af8;
  wire v85ac62;
  wire v872f22;
  wire v87622b;
  wire v87ed2d;
  wire v873227;
  wire v859a0a;
  wire v87313e;
  wire v872c10;
  wire v87ed0e;
  wire v87e83a;
  wire v8728b4;
  wire v87ec1d;
  wire v868ba6;
  wire v8733d5;
  wire v873228;
  wire v87e816;
  wire v852cab;
  wire v872e15;
  wire v87287d;
  wire v85ac98;
  wire v87ec2a;
  wire v87304a;
  wire v87ed9c;
  wire v86854e;
  wire v87ed58;
  wire v87ec03;
  wire v87ecac;
  wire v85ad2e;
  wire v87eee5;
  wire v87e8ce;
  wire v8737cc;
  wire v87ecb7;
  wire v856902;
  wire v856893;
  wire v87ec93;
  wire v87e8aa;
  wire v8737d4;
  wire v87295c;
  wire v87ece1;
  wire v873291;
  wire v852d8b;
  wire v872d0b;
  wire v87ecfc;
  wire v872964;
  wire v872c9f;
  wire v87ed68;
  wire v87ef15;
  wire v87edcf;
  wire v868ace;
  wire v8732c5;
  wire v873181;
  wire v87ed81;
  wire v868b13;
  wire v87291d;
  wire v87939c;
  wire v873342;
  wire v87eda8;
  wire v858363;
  wire v8598fe;
  wire v872c73;
  wire v87ed6c;
  wire v87ed2c;
  wire v8728f3;
  wire v872f14;
  wire v87ec08;
  wire v8731cd;
  wire v87ec55;
  wire v875270;
  wire v872de7;
  wire v868b88;
  wire v858cf2;
  wire v873238;
  wire v87ed55;
  wire v868be9;
  wire v874d66;
  wire v872d34;
  wire v87e7e0;
  wire v874226;
  wire v844f9e;
  wire v87323a;
  wire v87ef04;
  wire v852af2;
  wire v87ecbe;
  wire v87ed87;
  wire v87ed6a;
  wire v87ed22;
  wire v8731e2;
  wire v87edb8;
  wire v8727fb;
  wire v87edbb;
  wire v87ed89;
  wire v85a55b;
  wire v87df12;
  wire v8736d4;
  wire v854114;
  wire v873298;
  wire v868bcc;
  wire v85884d;
  wire v87ec97;
  wire v8728aa;
  wire v85b0b9;
  wire v87e811;
  wire v87ee53;
  wire v872863;
  wire v87ec70;
  wire v87ec04;
  wire v87ec5b;
  wire v87ec88;
  wire v87ec67;
  wire v87291c;
  wire v868b6a;
  wire v87ece4;
  wire v8731f5;
  wire v87e894;
  wire v874056;
  wire v868b76;
  wire v87ef41;
  wire v872836;
  wire v87ed6d;
  wire v87edbf;
  wire v87ec3a;
  wire v87293b;
  wire v87ed15;
  wire v868bc5;
  wire v852651;
  wire v844fa5;
  wire v844f95;
  wire v872d50;
  wire v852613;
  wire v853e70;
  wire v873169;
  wire v87332a;
  wire v876227;
  wire v87ec5c;
  wire v8731ae;
  wire v873383;
  wire v87ec60;
  wire v87292f;
  wire v873042;
  wire v87ef7a;
  wire v844f97;
  wire v87ec34;
  wire v87332c;
  wire v873319;
  wire v872915;
  wire v87ec82;
  wire v87eca9;
  wire v87ece6;
  wire v87ecb3;
  wire v87ef71;
  wire v85259e;
  wire v87ec3d;
  wire v87ee8e;
  wire v8793ad;
  wire v844fa7;
  wire v87ef46;
  wire v87ec0f;
  wire v872b6a;
  wire v87ec59;
  wire v873118;
  wire v872cd4;
  wire v872c3b;
  wire v87e920;
  wire v87ef9b;
  wire v8737a3;
  wire v87edd3;
  wire v857022;
  wire v872f59;
  wire v855880;
  wire v87304f;
  wire v868ac6;
  wire v872ddf;
  wire v872822;
  wire v87630b;
  wire v87e838;
  wire v87ef70;
  wire v87eca5;
  wire v8730d5;
  wire v872fc4;
  wire v872f06;
  wire v87ec63;
  wire v87ec22;
  wire v852632;
  wire v87ec20;
  wire v87eda1;
  wire v87df27;
  wire v87ece5;
  wire v874053;
  wire v87eca6;
  wire v872ea3;
  wire v857e91;
  wire v872c18;
  wire v8685f8;
  wire v87eea7;
  wire v872fb2;
  wire v868b41;
  wire v8732f1;
  wire v8525f0;
  wire v868bce;
  wire v872856;
  wire v87ed98;
  wire v874047;
  wire v872de2;
  wire v868b0e;
  wire v87ef9a;
  wire v87edae;
  wire v872873;
  wire v87e7f6;
  wire v8731e1;
  wire v874063;
  wire v87b3e9;
  wire v868bac;
  wire v8598ae;
  wire v855c5b;
  wire v87ed40;
  wire v873189;
  wire v8732cb;
  wire v87edb0;
  wire v8737e1;
  wire v87aed9;
  wire v844fa9;
  wire v87eeef;
  wire v872f1f;
  wire v87ee04;
  wire v87ec46;
  wire v87ecab;
  wire v8731cf;
  wire v87ed71;
  wire v87ee13;
  wire v858aae;
  wire v87ebf7;
  wire v872cf6;
  wire v873126;
  wire v872cdb;
  wire v875285;
  wire v87ecfe;
  wire v858c10;
  wire v8732c6;
  wire v87ecb2;
  wire v872f42;
  wire v87281e;
  wire v87ed95;
  wire v874c36;
  wire v87459e;
  wire v87e8f4;
  wire v87ebf3;
  wire v872830;
  wire v87ece0;
  wire v868aef;
  wire v8737d6;
  wire v87ed19;
  wire v8731e8;
  wire v87eeed;
  wire v873058;
  wire v87edd1;
  wire v87ec35;
  wire v872921;
  wire v87ebe8;
  wire v873746;
  wire v87ec50;
  wire v872f89;
  wire v87624a;
  reg StoB_REQ0_p;
  input StoB_REQ0_n;
  reg StoB_REQ1_p;
  input StoB_REQ1_n;
  reg StoB_REQ2_p;
  input StoB_REQ2_n;
  reg StoB_REQ3_p;
  input StoB_REQ3_n;
  reg RtoB_ACK0_p;
  input RtoB_ACK0_n;
  reg RtoB_ACK1_p;
  input RtoB_ACK1_n;
  reg FULL_p;
  input FULL_n;
  reg EMPTY_p;
  input EMPTY_n;
  reg BtoS_ACK0_p;
  output BtoS_ACK0_n;
  reg BtoS_ACK1_p;
  output BtoS_ACK1_n;
  reg BtoS_ACK2_p;
  output BtoS_ACK2_n;
  reg BtoS_ACK3_p;
  output BtoS_ACK3_n;
  reg BtoR_REQ0_p;
  output BtoR_REQ0_n;
  reg BtoR_REQ1_p;
  output BtoR_REQ1_n;
  reg stateG7_0_p;
  output stateG7_0_n;
  reg stateG7_1_p;
  output stateG7_1_n;
  reg ENQ_p;
  output ENQ_n;
  reg DEQ_p;
  output DEQ_n;
  reg stateG12_p;
  output stateG12_n;
  reg SLC0_p;
  output SLC0_n;
  reg SLC1_p;
  output SLC1_n;
  reg jx0_p;
  output jx0_n;
  reg jx1_p;
  output jx1_n;
  reg jx2_p;
  output jx2_n;
  wire SLC0_n;
  wire ENQ_n;
  wire SLC1_n;

assign v87ec88 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & !v87323a;
assign v87ef0a = StoB_REQ2_p & v85a673 | !StoB_REQ2_p & v87ec1c;
assign v87ed7a = StoB_REQ2_p & v868aba | !StoB_REQ2_p & v844f91;
assign v8757c5 = StoB_REQ0_p & v872e81 | !StoB_REQ0_p & v853052;
assign v874053 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v87ece5;
assign v855989 = StoB_REQ2_p & v873723 | !StoB_REQ2_p & v868ba1;
assign v87ef9c = StoB_REQ3_p & v856f49 | !StoB_REQ3_p & v87ec4a;
assign v87e811 = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v85b0b9;
assign v87ebf7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v858aae;
assign v87edd5 = BtoS_ACK0_p & v87289c | !BtoS_ACK0_p & v873392;
assign v87304a = BtoS_ACK0_p & v87e86b | !BtoS_ACK0_p & v87ec2a;
assign BtoR_REQ1_n = !v852651;
assign v872878 = jx0_p & v844f91 | !jx0_p & v872d99;
assign v87e838 = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v87ec34;
assign v873250 = StoB_REQ0_p & v868aba | !StoB_REQ0_p & v8736f8;
assign v852651 = jx2_p & v85ac98 | !jx2_p & v868bc5;
assign v858bae = BtoS_ACK1_p & v87ec12 | !BtoS_ACK1_p & v8733af;
assign v87ecfc = jx0_p & v872d0b | !jx0_p & v87ebf6;
assign v873327 = StoB_REQ2_p & v852d87 | !StoB_REQ2_p & v8733e9;
assign v872fe0 = StoB_REQ0_p & v87ef83 | !StoB_REQ0_p & v872eb0;
assign v844fad = BtoR_REQ0_p & v844f91 | !BtoR_REQ0_p & !v844f91;
assign BtoS_ACK2_n = !v876322;
assign v844f9d = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v844f91;
assign v87ed83 = StoB_REQ1_p & v8588f4 | !StoB_REQ1_p & v87ecd1;
assign v874063 = ENQ_p & v8685f8 | !ENQ_p & v8731e1;
assign v87e894 = BtoS_ACK0_p & v87ec5b | !BtoS_ACK0_p & !v8731f5;
assign v87289c = StoB_REQ1_p & v87302a | !StoB_REQ1_p & v8757ca;
assign v8525f0 = StoB_REQ1_p & v8733da | !StoB_REQ1_p & v872837;
assign v87287d = DEQ_p & v87313e | !DEQ_p & v872e15;
assign v87edcf = BtoS_ACK3_p & v8752ab | !BtoS_ACK3_p & v868aba;
assign v858bc4 = BtoS_ACK1_p & v87ecd1 | !BtoS_ACK1_p & v87ec53;
assign v87ed9e = StoB_REQ1_p & v87edd0 | !StoB_REQ1_p & v87eec0;
assign v87eee0 = StoB_REQ0_p & v872d64 | !StoB_REQ0_p & v8737e3;
assign v87939c = BtoS_ACK2_p & v87eeaa | !BtoS_ACK2_p & v87e86b;
assign v87295c = BtoS_ACK0_p & v868aba | !BtoS_ACK0_p & v8737d4;
assign v8732f1 = jx0_p & v87ed61 | !jx0_p & !v868b41;
assign v872ec9 = BtoS_ACK1_p & v852d87 | !BtoS_ACK1_p & v87ec0a;
assign v87ed3e = StoB_REQ0_p & v873799 | !StoB_REQ0_p & v8736f4;
assign v87ed04 = jx0_p & v87ed61 | !jx0_p & v844f91;
assign v872bf1 = BtoS_ACK0_p & v87ed9e | !BtoS_ACK0_p & v85724c;
assign v872e0f = BtoS_ACK0_p & v872d64 | !BtoS_ACK0_p & v872fa1;
assign v852226 = StoB_REQ1_p & v87ec2d | !StoB_REQ1_p & v87ed80;
assign v87ec32 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8733da;
assign v844fb3 = stateG7_1_p & v844f91 | !stateG7_1_p & !v844f91;
assign v87ecbf = BtoS_ACK1_p & v872fa7 | !BtoS_ACK1_p & v8728a3;
assign v87ed75 = BtoS_ACK0_p & v85b5e0 | !BtoS_ACK0_p & v87622d;
assign v844f91 = 1;
assign v87630b = DEQ_p & v872ddf | !DEQ_p & v872822;
assign v87ec8e = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v873779;
assign v87eeed = EMPTY_p & v8737d6 | !EMPTY_p & !v8731e8;
assign v873383 = StoB_REQ0_p & v844f99 | !StoB_REQ0_p & v844f91;
assign v87ec1a = StoB_REQ1_p & v87ed5b | !StoB_REQ1_p & v852d6f;
assign v87305a = BtoS_ACK1_p & v872d64 | !BtoS_ACK1_p & v87e8e1;
assign v872e15 = EMPTY_p & v859a0a | !EMPTY_p & !v852cab;
assign v87332f = BtoS_ACK1_p & v87ec98 | !BtoS_ACK1_p & v872d03;
assign v87ebe4 = StoB_REQ3_p & v87338a | !StoB_REQ3_p & v872c60;
assign v85b091 = StoB_REQ2_p & v87ed48 | !StoB_REQ2_p & v852d87;
assign v872e6f = StoB_REQ3_p & v856f49 | !StoB_REQ3_p & v874242;
assign v874c36 = DEQ_p & v87281e | !DEQ_p & v87ed95;
assign v87283c = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844f9f;
assign v8731e1 = jx1_p & v868b0e | !jx1_p & v87e7f6;
assign v87ec23 = StoB_REQ1_p & v87ed1c | !StoB_REQ1_p & v87322c;
assign v87eee6 = EMPTY_p & v844f91 | !EMPTY_p & !v844fb9;
assign v868adc = jx0_p & v852d67 | !jx0_p & v87ed96;
assign v87332a = DEQ_p & v872d50 | !DEQ_p & v873169;
assign v87ec59 = stateG12_p & v87ef46 | !stateG12_p & !v872b6a;
assign v876245 = BtoS_ACK1_p & v87ed5b | !BtoS_ACK1_p & v872e81;
assign v87ed10 = BtoS_ACK0_p & v87edf9 | !BtoS_ACK0_p & v87ec06;
assign v87ec4a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v8752ab;
assign v874c37 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v87ed3e;
assign v87ec12 = StoB_REQ2_p & v872c60 | !StoB_REQ2_p & v87ecd7;
assign v8732c6 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v873071;
assign v87ed55 = StoB_REQ2_p & v87ed9f | !StoB_REQ2_p & v844f91;
assign v853eb8 = StoB_REQ0_p & v868b30 | !StoB_REQ0_p & v85a712;
assign v868b88 = BtoS_ACK1_p & v8728f3 | !BtoS_ACK1_p & v872de7;
assign v872ee9 = jx0_p & v872f13 | !jx0_p & v872d64;
assign v873118 = DEQ_p & v87ec59 | !DEQ_p & v87ef46;
assign v87ece1 = StoB_REQ0_p & v87eeaa | !StoB_REQ0_p & v873176;
assign v87ee02 = BtoS_ACK3_p & v8752ab | !BtoS_ACK3_p & !v872c60;
assign v87efcc = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v873250;
assign v873078 = EMPTY_p & v87edc6 | !EMPTY_p & v872d64;
assign v87ec63 = jx0_p & v872f06 | !jx0_p & v844f91;
assign v87ec0f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87ec34;
assign v87ebef = BtoS_ACK1_p & v87302a | !BtoS_ACK1_p & v852227;
assign v8686b4 = jx1_p & v87eccf | !jx1_p & v8728c0;
assign v8731d4 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v872c60;
assign v872c60 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87ec9f;
assign BtoS_ACK3_n = !v87624a;
assign v87307b = StoB_REQ3_p & v8745a5 | !StoB_REQ3_p & v8733e9;
assign v8745a9 = StoB_REQ1_p & v872c60 | !StoB_REQ1_p & v872f69;
assign v87ec04 = jx0_p & v87ec70 | !jx0_p & v859a0a;
assign v87ed6d = FULL_p & v87e83a | !FULL_p & v872836;
assign v8733d5 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v868ba6;
assign v872ecb = StoB_REQ1_p & v856f49 | !StoB_REQ1_p & v8732f0;
assign v87323e = BtoS_ACK0_p & v87ed83 | !BtoS_ACK0_p & v856718;
assign v844fa5 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f91;
assign v8750ad = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & v844fab;
assign v872d4f = stateG7_1_p & v876314 | !stateG7_1_p & v844f9f;
assign v857beb = StoB_REQ2_p & v87338a | !StoB_REQ2_p & !v868aba;
assign v872877 = stateG12_p & v874c38 | !stateG12_p & v8757d7;
assign v872cf6 = StoB_REQ0_p & v87eeef | !StoB_REQ0_p & v87ebf7;
assign v8752b0 = BtoS_ACK1_p & v872fa7 | !BtoS_ACK1_p & v874bf2;
assign v873746 = DEQ_p & v87ed71 | !DEQ_p & v87ebe8;
assign v873042 = EMPTY_p & v87292f | !EMPTY_p & v844f91;
assign v87ec95 = jx0_p & v87ec14 | !jx0_p & v8757d2;
assign v873058 = DEQ_p & v87ebf3 | !DEQ_p & v87eeed;
assign v87ed5b = StoB_REQ3_p & v87338a | !StoB_REQ3_p & v872e81;
assign v872e9a = BtoS_ACK1_p & v87ed62 | !BtoS_ACK1_p & v872c81;
assign v872ff7 = BtoS_ACK0_p & v872f79 | !BtoS_ACK0_p & v873176;
assign v868b71 = StoB_REQ0_p & v872d67 | !StoB_REQ0_p & v8730b0;
assign v8731f8 = StoB_REQ2_p & v856f49 | !StoB_REQ2_p & v8728cb;
assign v87ee84 = StoB_REQ3_p & v87378d | !StoB_REQ3_p & v844f91;
assign v844f9e = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & !v844f91;
assign v872cdb = DEQ_p & v87ee13 | !DEQ_p & v873126;
assign v872f82 = BtoS_ACK2_p & v87ebf5 | !BtoS_ACK2_p & v8588f4;
assign v86854e = BtoS_ACK0_p & v872f79 | !BtoS_ACK0_p & v87ed9c;
assign v857e91 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v87ec34;
assign v87ec5b = StoB_REQ1_p & v87323a | !StoB_REQ1_p & !v873375;
assign v87422b = jx0_p & v855c35 | !jx0_p & v872c17;
assign v844fb9 = stateG12_p & v844f91 | !stateG12_p & !v844f91;
assign v8728a3 = StoB_REQ1_p & v872e81 | !StoB_REQ1_p & v87eddd;
assign v87eeaa = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & v872fb8;
assign v87ed70 = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & v87291a;
assign v87ed3f = BtoS_ACK2_p & v873327 | !BtoS_ACK2_p & v87e8f3;
assign v8728f3 = StoB_REQ2_p & v87ed2c | !StoB_REQ2_p & v8538fd;
assign v8731e8 = jx0_p & v87ed19 | !jx0_p & v844f91;
assign v87edd3 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v8737a3;
assign v872936 = EMPTY_p & v8731fb | !EMPTY_p & v87ed04;
assign v87ed87 = BtoS_ACK1_p & v852af2 | !BtoS_ACK1_p & v87ecbe;
assign v87ecb1 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87ed70;
assign v85b2d3 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8730eb;
assign v868b3d = StoB_REQ2_p & v8564be | !StoB_REQ2_p & v873726;
assign v857ea2 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v85271e;
assign v858c10 = ENQ_p & v872cdb | !ENQ_p & v87ecfe;
assign v8728d6 = jx0_p & v872ec1 | !jx0_p & v872fa5;
assign v873379 = StoB_REQ3_p & v87eeaa | !StoB_REQ3_p & v868aba;
assign v8737c6 = StoB_REQ2_p & v856f49 | !StoB_REQ2_p & v87307b;
assign v87eca2 = BtoS_ACK2_p & v8730c6 | !BtoS_ACK2_p & v85b091;
assign v87ed8f = EMPTY_p & v8757d7 | !EMPTY_p & v872877;
assign v87ec50 = jx1_p & v873058 | !jx1_p & !v873746;
assign v868bc5 = ENQ_p & v872c9f | !ENQ_p & v87ed15;
assign v872e8e = ENQ_p & v8686b4 | !ENQ_p & v87ed23;
assign v87287b = BtoS_ACK2_p & v87eccb | !BtoS_ACK2_p & v87ed13;
assign v856893 = jx0_p & v87e8ce | !jx0_p & v856902;
assign v87ecef = BtoS_ACK2_p & v854111 | !BtoS_ACK2_p & v87ed3d;
assign v87ec89 = stateG7_1_p & v844faf | !stateG7_1_p & v87eca1;
assign v844f99 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f91;
assign v873126 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v872cf6;
assign v868be9 = BtoS_ACK1_p & v87ed55 | !BtoS_ACK1_p & v868af8;
assign v8736f4 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v868b29;
assign v873392 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v853052;
assign v8564be = StoB_REQ3_p & v87302a | !StoB_REQ3_p & v8757c6;
assign v87ecfd = StoB_REQ0_p & v87332f | !StoB_REQ0_p & v853052;
assign v87ef70 = jx0_p & v87e838 | !jx0_p & v872b6a;
assign v85259e = DEQ_p & v872915 | !DEQ_p & v87ef71;
assign v87edcc = BtoS_ACK0_p & v872ee2 | !BtoS_ACK0_p & v872da9;
assign v868b30 = BtoS_ACK1_p & v872e81 | !BtoS_ACK1_p & v852227;
assign v852632 = DEQ_p & v87ef70 | !DEQ_p & v87ec22;
assign v87ec2c = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & !v86e02d;
assign v8732f0 = BtoS_ACK2_p & v8745a5 | !BtoS_ACK2_p & v87ed3d;
assign v87eec0 = StoB_REQ2_p & v87ec98 | !StoB_REQ2_p & v852d87;
assign v87ed84 = BtoS_ACK1_p & v872e81 | !BtoS_ACK1_p & v87ed2f;
assign v859412 = BtoS_ACK2_p & v872f67 | !BtoS_ACK2_p & v8731f8;
assign v87e8be = StoB_REQ0_p & v8731c8 | !StoB_REQ0_p & v872f17;
assign v872e22 = StoB_REQ1_p & v87302a | !StoB_REQ1_p & v872e81;
assign v87ee53 = jx0_p & v87e811 | !jx0_p & v859a0a;
assign v87ebf6 = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & v87ec8e;
assign v873291 = BtoS_ACK0_p & v872f79 | !BtoS_ACK0_p & v87ece1;
assign v872de7 = StoB_REQ1_p & v87ec55 | !StoB_REQ1_p & v87bbdd;
assign v87eda8 = BtoS_ACK1_p & v87bbdd | !BtoS_ACK1_p & v873342;
assign v8731cd = StoB_REQ2_p & v87eeaa | !StoB_REQ2_p & v87ec08;
assign v87623a = StoB_REQ1_p & v87ed62 | !StoB_REQ1_p & v87ec12;
assign v87eccf = DEQ_p & v8728d6 | !DEQ_p & v87422b;
assign v87500a = StoB_REQ1_p & v873333 | !StoB_REQ1_p & v87ed97;
assign v859947 = StoB_REQ2_p & v844f9b | !StoB_REQ2_p & v844f91;
assign v87ebee = RtoB_ACK0_n & v844f9f | !RtoB_ACK0_n & v87ed79;
assign v868b92 = DEQ_p & v8582c0 | !DEQ_p & v872dd8;
assign v87e83a = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & v87ed0e;
assign v87ecab = BtoS_ACK1_p & v87ee04 | !BtoS_ACK1_p & v87ec46;
assign v87e855 = StoB_REQ2_p & v856f49 | !StoB_REQ2_p & v8733e9;
assign v87ec42 = BtoS_ACK0_p & v872fa7 | !BtoS_ACK0_p & v853eb8;
assign v85a0a4 = stateG7_0_p & v844fb3 | !stateG7_0_p & v844f91;
assign v853052 = BtoS_ACK1_p & v872fa7 | !BtoS_ACK1_p & v8732c4;
assign v85b0b9 = StoB_REQ0_p & v8728aa | !StoB_REQ0_p & v87ed2d;
assign v87ec53 = StoB_REQ1_p & v872f82 | !StoB_REQ1_p & v87ec6d;
assign v87ec6d = BtoS_ACK2_p & v872975 | !BtoS_ACK2_p & v87ecd1;
assign v856719 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v872c19;
assign BtoS_ACK0_n = v8793ad;
assign v87292f = jx0_p & v8731ae | !jx0_p & v87ec60;
assign v868ae0 = jx0_p & v868b4a | !jx0_p & v8730c8;
assign v872ddf = jx0_p & v857022 | !jx0_p & v868ac6;
assign v8733e9 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v875111;
assign v872f06 = FULL_p & v872fc4 | !FULL_p & !v87e838;
assign v87ec93 = DEQ_p & v87ed58 | !DEQ_p & !v856893;
assign v85448e = BtoS_ACK1_p & v8598e6 | !BtoS_ACK1_p & v87efce;
assign v872ec1 = BtoS_ACK0_p & v87eda9 | !BtoS_ACK0_p & v87ebfe;
assign v85ad2e = BtoS_ACK1_p & v873375 | !BtoS_ACK1_p & v87ecac;
assign v87302a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v87efc2;
assign v87eef6 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f99;
assign v873293 = StoB_REQ2_p & v8750ad | !StoB_REQ2_p & v844f9b;
assign v8733af = StoB_REQ1_p & v872c60 | !StoB_REQ1_p & v87ed51;
assign v852613 = stateG12_p & v844fa5 | !stateG12_p & !v872d50;
assign v872c51 = BtoS_ACK1_p & v87edd0 | !BtoS_ACK1_p & v872dff;
assign v87ed95 = jx0_p & v873126 | !jx0_p & v87ecb2;
assign v87ed98 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v872856;
assign v868bce = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8525f0;
assign v87ec06 = StoB_REQ0_p & v872890 | !StoB_REQ0_p & v872e7a;
assign v87eca1 = BtoR_REQ1_p & v844f9f | !BtoR_REQ1_p & !v844f91;
assign v873375 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v872d35;
assign v87e8aa = StoB_REQ1_p & v87eeaa | !StoB_REQ1_p & v868bde;
assign v87ed06 = EMPTY_p & v844f91 | !EMPTY_p & v872d64;
assign v87313e = stateG12_p & v859a0a | !stateG12_p & v87efcc;
assign v87ecbd = BtoS_ACK3_p & v86e02d | !BtoS_ACK3_p & v8733e9;
assign v87624a = jx2_p & v858c10 | !jx2_p & v872f89;
assign v87ec5c = StoB_REQ0_p & v844f9b | !StoB_REQ0_p & v844f91;
assign v87ed9c = BtoS_ACK1_p & v868aba | !BtoS_ACK1_p & v868bde;
assign v87ed61 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v87ec32;
assign v855c5b = jx0_p & v87ed98 | !jx0_p & v844f91;
assign v85b574 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v8733ec;
assign v872f4c = StoB_REQ1_p & v87ec98 | !StoB_REQ1_p & v872fa7;
assign v85b5e0 = StoB_REQ1_p & v8733e9 | !StoB_REQ1_p & v879395;
assign v872f17 = BtoS_ACK1_p & v87ed76 | !BtoS_ACK1_p & v87ed9d;
assign v873228 = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & v8733d5;
assign v872856 = StoB_REQ0_p & v87ec32 | !StoB_REQ0_p & v868bce;
assign v8737d4 = BtoS_ACK1_p & v872f79 | !BtoS_ACK1_p & v87e8aa;
assign v8732d3 = stateG7_0_p & v85409b | !stateG7_0_p & v852e67;
assign v87323a = RtoB_ACK0_p & v844f9e | !RtoB_ACK0_p & v87eeaa;
assign v8737c4 = jx0_p & v872d56 | !jx0_p & v844f91;
assign v872d7f = StoB_REQ2_p & v87ee8b | !StoB_REQ2_p & v872ed3;
assign v87ecdb = StoB_REQ1_p & v87eda6 | !StoB_REQ1_p & v87ed45;
assign v874056 = FULL_p & v87e83a | !FULL_p & !v87e894;
assign v872fee = StoB_REQ0_p & v87ed84 | !StoB_REQ0_p & v872ec9;
assign v8732cb = jx0_p & v87edae | !jx0_p & v844f91;
assign v872d99 = FULL_p & v87edc4 | !FULL_p & !v844f99;
assign v872f59 = StoB_REQ1_p & v844f99 | !StoB_REQ1_p & v844f91;
assign v87ebe8 = EMPTY_p & v872921 | !EMPTY_p & v844f91;
assign v87338a = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v87eeaa;
assign v87eda4 = BtoS_ACK0_p & v87eef6 | !BtoS_ACK0_p & v85b574;
assign v87e8f3 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v8733e9;
assign v8750bd = DEQ_p & v844f91 | !DEQ_p & v87ed06;
assign v8737cc = BtoS_ACK1_p & v872d35 | !BtoS_ACK1_p & v8732c2;
assign v844fa7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f91;
assign v85abe7 = stateG7_1_p & v876314 | !stateG7_1_p & v844f91;
assign v87ec11 = BtoS_ACK0_p & v87289c | !BtoS_ACK0_p & v87ecfd;
assign v8737e1 = ENQ_p & v8598ae | !ENQ_p & v87edb0;
assign v85ab45 = StoB_REQ3_p & v87302a | !StoB_REQ3_p & v857ea2;
assign v873799 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & v8750ad;
assign v87ecb7 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v8737cc;
assign v87ed6b = BtoS_ACK2_p & v87ed3b | !BtoS_ACK2_p & v87ed7a;
assign v87ecc3 = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v872fa7;
assign v87ebf5 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v87302a;
assign v87ee9d = StoB_REQ2_p & v857ea2 | !StoB_REQ2_p & v872ed3;
assign v8752ab = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & v85a0a4;
assign v8731b2 = DEQ_p & v87ed01 | !DEQ_p & v872936;
assign v87e8d0 = BtoS_ACK0_p & v87ec1a | !BtoS_ACK0_p & v872f5d;
assign v87ed7b = StoB_REQ0_p & v876245 | !StoB_REQ0_p & v87ec6b;
assign v879395 = StoB_REQ2_p & v8733e9 | !StoB_REQ2_p & v87ed27;
assign v87379c = BtoS_ACK2_p & v8733e9 | !BtoS_ACK2_p & v87ec05;
assign v8731c8 = BtoS_ACK1_p & v868b8b | !BtoS_ACK1_p & v872e6f;
assign v87330a = jx1_p & v8737c4 | !jx1_p & v844f91;
assign v87e7e0 = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v872d34;
assign v844faf = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & !v844f91;
assign v872df4 = jx1_p & v87ec49 | !jx1_p & v873784;
assign v872c81 = BtoS_ACK2_p & v872c60 | !BtoS_ACK2_p & v87ed62;
assign v872fa5 = BtoS_ACK0_p & v87ed62 | !BtoS_ACK0_p & v87e85d;
assign v873189 = DEQ_p & v87ed04 | !DEQ_p & v87ed40;
assign v87edb2 = DEQ_p & v87eccc | !DEQ_p & v8757d4;
assign v876322 = jx2_p & v87377f | !jx2_p & v87372e;
assign v87efce = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v87eceb;
assign v87eee5 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v85ad2e;
assign v87622b = StoB_REQ1_p & v868af8 | !StoB_REQ1_p & v872f22;
assign v8582c0 = stateG12_p & v872dd8 | !stateG12_p & v87eda4;
assign v872873 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v844f95;
assign v872d50 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844f95;
assign v87ece4 = BtoS_ACK1_p & v873375 | !BtoS_ACK1_p & v868b6a;
assign v87edcb = stateG7_0_p & v844fb3 | !stateG7_0_p & !v844fb3;
assign v872c18 = jx0_p & v857e91 | !jx0_p & !v872d50;
assign v872cd6 = StoB_REQ1_p & v872e81 | !StoB_REQ1_p & v87379c;
assign v872b6a = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & !v87ec0f;
assign v87ec6b = BtoS_ACK1_p & v852d6f | !BtoS_ACK1_p & v872cd6;
assign v87ecd1 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v852d87;
assign v85271e = stateG7_0_p & v85abe7 | !stateG7_0_p & v872d4f;
assign v87ed6c = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v8752ab;
assign v872975 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v85ab45;
assign v8727f7 = StoB_REQ0_p & v872e81 | !StoB_REQ0_p & v87ecbf;
assign v87eca9 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v87ec82;
assign v87291f = BtoS_ACK0_p & v87ecfa | !BtoS_ACK0_p & v873177;
assign v872f67 = StoB_REQ2_p & v856f49 | !StoB_REQ2_p & v857ea2;
assign v86e02d = stateG7_0_p & v873197 | !stateG7_0_p & v872f4e;
assign v872f1a = EMPTY_p & v87ed75 | !EMPTY_p & v87e8f1;
assign v87bbdd = StoB_REQ2_p & v868aba | !StoB_REQ2_p & v8538fd;
assign v87ed19 = FULL_p & v873172 | !FULL_p & !v844f9b;
assign v87ec51 = stateG12_p & v872b5c | !stateG12_p & v87ec72;
assign v87ec5a = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v8598e6;
assign v872e7a = BtoS_ACK1_p & v87ee9d | !BtoS_ACK1_p & v8733c1;
assign v87ed68 = BtoS_ACK2_p & v87e86b | !BtoS_ACK2_p & v872f79;
assign BtoR_REQ0_n = !v868bef;
assign v8731f5 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v87ece4;
assign v87372a = BtoS_ACK1_p & v852d6f | !BtoS_ACK1_p & v87ec23;
assign v868b13 = StoB_REQ0_p & v87ef15 | !StoB_REQ0_p & v87ed81;
assign v8727fb = StoB_REQ1_p & v87338a | !StoB_REQ1_p & !v87edb8;
assign v868ba6 = BtoS_ACK1_p & v873375 | !BtoS_ACK1_p & v87ec1d;
assign v872de4 = StoB_REQ3_p & v87ec2d | !StoB_REQ3_p & v872c60;
assign v87ecfa = StoB_REQ1_p & v85a673 | !StoB_REQ1_p & v87ef0a;
assign v87ec19 = StoB_REQ3_p & v87ec2d | !StoB_REQ3_p & !v87ee02;
assign v873077 = StoB_REQ2_p & v87ec19 | !StoB_REQ2_p & v87ecd7;
assign v868b6a = StoB_REQ1_p & v87291c | !StoB_REQ1_p & v873375;
assign v8737e4 = StoB_REQ2_p & v8564be | !StoB_REQ2_p & v85a673;
assign v85ac62 = BtoS_ACK1_p & v868aba | !BtoS_ACK1_p & v868af8;
assign v87ec65 = StoB_REQ1_p & v868aba | !StoB_REQ1_p & v87bbdd;
assign v8730c8 = FULL_p & v87323e | !FULL_p & v872bf1;
assign v872db6 = StoB_REQ2_p & v87307b | !StoB_REQ2_p & v87ed27;
assign v873741 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v85adeb;
assign v87291c = BtoS_ACK2_p & v87ec88 | !BtoS_ACK2_p & v87ec67;
assign v872b76 = jx2_p & v879392 | !jx2_p & !v87ecde;
assign v873759 = BtoS_ACK1_p & v857ea2 | !BtoS_ACK1_p & v859412;
assign v87edd7 = BtoS_ACK1_p & v87ec12 | !BtoS_ACK1_p & v8745a9;
assign v87ed71 = BtoS_ACK0_p & v87ec46 | !BtoS_ACK0_p & v8731cf;
assign v872836 = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & !v87ef41;
assign v873181 = StoB_REQ1_p & v87ed68 | !StoB_REQ1_p & v8732c5;
assign v872f22 = StoB_REQ2_p & v873379 | !StoB_REQ2_p & v8538fd;
assign v8728cb = StoB_REQ3_p & v856f49 | !StoB_REQ3_p & v857ea2;
assign v87edbb = StoB_REQ3_p & v87338a | !StoB_REQ3_p & !v87323a;
assign v87ecb2 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v8732c6;
assign v87eca5 = StoB_REQ1_p & v872d64 | !StoB_REQ1_p & v844f91;
assign v87ec34 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v844f97;
assign v844f9f = RtoB_ACK1_p & v844f91 | !RtoB_ACK1_p & !v844f91;
assign v868b76 = BtoS_ACK1_p & v87323a | !BtoS_ACK1_p & !v87291c;
assign v874bf2 = StoB_REQ1_p & v872e81 | !StoB_REQ1_p & v876307;
assign v87ed3d = StoB_REQ2_p & v8745a5 | !StoB_REQ2_p & v87307b;
assign v87ecac = StoB_REQ1_p & v87338a | !StoB_REQ1_p & !v87ec03;
assign v8598fe = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v858363;
assign v87286f = StoB_REQ3_p & v87ecb1 | !StoB_REQ3_p & v844f91;
assign v87ee13 = stateG12_p & v872f1f | !stateG12_p & v87ed71;
assign v872e8b = StoB_REQ2_p & v873723 | !StoB_REQ2_p & v87ed5b;
assign v872c9f = jx1_p & v87ec93 | !jx1_p & v872964;
assign v87ed0e = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v872c10;
assign v8737ab = StoB_REQ1_p & v872dff | !StoB_REQ1_p & v87eca2;
assign v852d8b = jx0_p & v87295c | !jx0_p & v873291;
assign v87ed23 = jx1_p & v8594bd | !jx1_p & v8525dc;
assign v87aed9 = jx2_p & v844f91 | !jx2_p & !v8737e1;
assign v87df27 = jx2_p & v87e920 | !jx2_p & v87eda1;
assign v87ec25 = StoB_REQ1_p & v868b8b | !StoB_REQ1_p & v87ed76;
assign v874064 = DEQ_p & v87ec01 | !DEQ_p & !v87ebf6;
assign v87e816 = stateG12_p & v87e83a | !stateG12_p & v873228;
assign v87e8f1 = FULL_p & v876238 | !FULL_p & v872f60;
assign v872964 = DEQ_p & v852d8b | !DEQ_p & !v87ecfc;
assign v873227 = StoB_REQ0_p & v85ac62 | !StoB_REQ0_p & v87ed2d;
assign v872dd8 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v87eca7;
assign v87ece5 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f99;
assign v87622d = StoB_REQ0_p & v87ecd2 | !StoB_REQ0_p & v87ec0b;
assign v87ed6a = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v87ed87;
assign v87ef77 = StoB_REQ1_p & v87ed92 | !StoB_REQ1_p & v872f69;
assign v872c3b = DEQ_p & v872b6a | !DEQ_p & v872cd4;
assign v87efc9 = stateG7_1_p & v873370 | !stateG7_1_p & v844f91;
assign v8733da = BtoS_ACK2_p & v873293 | !BtoS_ACK2_p & v8750ad;
assign v87ec9f = RtoB_ACK0_n & v844f9f | !RtoB_ACK0_n & v8732d3;
assign v87e8e1 = StoB_REQ1_p & v872d64 | !StoB_REQ1_p & v87ecda;
assign v857f15 = BtoS_ACK1_p & v87ec2d | !BtoS_ACK1_p & v852226;
assign v85ac98 = ENQ_p & v874064 | !ENQ_p & v87287d;
assign v87ede2 = BtoS_ACK1_p & v859947 | !BtoS_ACK1_p & v872ee2;
assign v856902 = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & v87ecb7;
assign v87ed58 = jx0_p & v87304a | !jx0_p & v86854e;
assign v8728b4 = BtoS_ACK2_p & v873375 | !BtoS_ACK2_p & v857beb;
assign v87efc2 = stateG7_0_p & v855cab | !stateG7_0_p & v87efc9;
assign v87ec05 = StoB_REQ2_p & v872e81 | !StoB_REQ2_p & v8733e9;
assign v874c38 = BtoS_ACK0_p & v87ec5a | !BtoS_ACK0_p & v873079;
assign v85a55b = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v87ed89;
assign v872fb2 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v87eea7;
assign v87eea7 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & v844f99;
assign v87e920 = ENQ_p & v873118 | !ENQ_p & !v872c3b;
assign v8731a1 = BtoS_ACK0_p & v87ed1e | !BtoS_ACK0_p & v87ec40;
assign v872890 = BtoS_ACK1_p & v856f49 | !BtoS_ACK1_p & v872ecb;
assign v87ec03 = BtoS_ACK2_p & v868aba | !BtoS_ACK2_p & !v857beb;
assign v852d93 = BtoS_ACK0_p & v87623a | !BtoS_ACK0_p & v872c93;
assign v8731e2 = FULL_p & v87e83a | !FULL_p & v87ed22;
assign DEQ_n = !v862858;
assign v87ecd7 = StoB_REQ3_p & v872c60 | !StoB_REQ3_p & v844f91;
assign v873370 = BtoR_REQ1_p & v844f9f | !BtoR_REQ1_p & v844f91;
assign v85884d = EMPTY_p & v874226 | !EMPTY_p & !v868bcc;
assign v872921 = jx0_p & v87ec35 | !jx0_p & v87ed71;
assign v87ec20 = jx1_p & v87630b | !jx1_p & !v852632;
assign v87edb8 = StoB_REQ2_p & v87323a | !StoB_REQ2_p & !v872d35;
assign v87ec55 = BtoS_ACK2_p & v8731cd | !BtoS_ACK2_p & v872f79;
assign v872ea3 = jx0_p & v872d56 | !jx0_p & !v87eca6;
assign v868bcc = jx0_p & v8731e2 | !jx0_p & v873298;
assign v8589e8 = DEQ_p & v8728e2 | !DEQ_p & v872f1a;
assign v87ed36 = jx1_p & v8731b2 | !jx1_p & v844f91;
assign v872f1f = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v87eeef;
assign v872915 = jx0_p & v873319 | !jx0_p & v872d50;
assign v868baa = EMPTY_p & v872ee9 | !EMPTY_p & v872d64;
assign v86284b = BtoS_ACK0_p & v8732c4 | !BtoS_ACK0_p & v868af3;
assign v87eccb = StoB_REQ2_p & v8728cb | !StoB_REQ2_p & v872ed3;
assign v873774 = DEQ_p & v87eda4 | !DEQ_p & v87ecd5;
assign v85adeb = StoB_REQ0_p & v873799 | !StoB_REQ0_p & v85b2d3;
assign v87ec28 = DEQ_p & v87ec51 | !DEQ_p & v87ed8f;
assign v855880 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v872f59;
assign v87293b = DEQ_p & v87ee53 | !DEQ_p & v87ec3a;
assign v872c19 = BtoS_ACK1_p & v8598e6 | !BtoS_ACK1_p & v87ec5a;
assign v8730d5 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v87eca5;
assign v87ec2d = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v87ed9f;
assign v87ecea = StoB_REQ2_p & v872d64 | !StoB_REQ2_p & v873172;
assign v87ebfe = BtoS_ACK1_p & v87eda9 | !BtoS_ACK1_p & v872c81;
assign v8730f3 = StoB_REQ2_p & v87302a | !StoB_REQ2_p & v87ed48;
assign v87ecb5 = StoB_REQ1_p & v872d03 | !StoB_REQ1_p & v872fa7;
assign v87ef9b = StoB_REQ1_p & v844f9b | !StoB_REQ1_p & v844f91;
assign v87e85b = BtoS_ACK1_p & v87ef0a | !BtoS_ACK1_p & v87500a;
assign v87ed96 = FULL_p & v87edd5 | !FULL_p & v87ec11;
assign v873176 = BtoS_ACK1_p & v872f79 | !BtoS_ACK1_p & v868bde;
assign v873071 = BtoS_ACK2_p & v844f99 | !BtoS_ACK2_p & !v844f91;
assign v872e7f = BtoS_ACK1_p & v8588f4 | !BtoS_ACK1_p & v872f82;
assign v87eccc = jx0_p & v87edcc | !jx0_p & !v844f99;
assign v87ed62 = StoB_REQ2_p & v87ec2d | !StoB_REQ2_p & v872c60;
assign v87ebf4 = BtoS_ACK1_p & v87ed62 | !BtoS_ACK1_p & v852626;
assign v872e99 = StoB_REQ1_p & v872de4 | !StoB_REQ1_p & v872f69;
assign v87318f = BtoS_ACK1_p & v8757ca | !BtoS_ACK1_p & v87ecc3;
assign v87eca6 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & !v874053;
assign v87ec41 = StoB_REQ2_p & v86e02d | !StoB_REQ2_p & v844f9d;
assign v8728e2 = stateG12_p & v8567f5 | !stateG12_p & v87ec72;
assign v868ace = StoB_REQ3_p & v87eeaa | !StoB_REQ3_p & v87edcf;
assign v856f49 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v86e02d;
assign v87ed0b = StoB_REQ1_p & v8733e9 | !StoB_REQ1_p & v872db6;
assign v873784 = DEQ_p & v844f91 | !DEQ_p & v868baa;
assign v858cf2 = StoB_REQ0_p & v875270 | !StoB_REQ0_p & v868b88;
assign v8737e3 = BtoS_ACK1_p & v873172 | !BtoS_ACK1_p & v872d64;
assign v868bde = BtoS_ACK2_p & v868aba | !BtoS_ACK2_p & v872f79;
assign v87ed22 = BtoS_ACK0_p & v87ecbe | !BtoS_ACK0_p & v87ed6a;
assign v87ec96 = StoB_REQ2_p & v87ebe4 | !StoB_REQ2_p & v872c60;
assign v8731cf = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87ecab;
assign v844fa9 = BtoS_ACK2_p & v844f91 | !BtoS_ACK2_p & !v844f91;
assign v87ecda = BtoS_ACK2_p & v87ec1b | !BtoS_ACK2_p & v872d64;
assign v87ec49 = DEQ_p & v844f91 | !DEQ_p & v873078;
assign v872fa1 = StoB_REQ0_p & v872d64 | !StoB_REQ0_p & v87305a;
assign v87ef04 = StoB_REQ3_p & v87323a | !StoB_REQ3_p & v868aba;
assign v87edd0 = StoB_REQ2_p & v87302a | !StoB_REQ2_p & v872e81;
assign v85a673 = StoB_REQ3_p & v87302a | !StoB_REQ3_p & v872e81;
assign v87ec40 = StoB_REQ0_p & v857f15 | !StoB_REQ0_p & v87332b;
assign v87e7f6 = jx0_p & v87edae | !jx0_p & !v872873;
assign v873048 = BtoS_ACK1_p & v87ec12 | !BtoS_ACK1_p & v87ef77;
assign v8793a7 = StoB_REQ0_p & v87ebef | !StoB_REQ0_p & v87318f;
assign v872d67 = BtoS_ACK1_p & v872de4 | !BtoS_ACK1_p & v87eda9;
assign v8757d2 = BtoS_ACK0_p & v87ed62 | !BtoS_ACK0_p & v872e92;
assign v873197 = stateG7_1_p & v844faf | !stateG7_1_p & v844f91;
assign v87eda9 = StoB_REQ2_p & v87ec2d | !StoB_REQ2_p & v872de4;
assign v87ed89 = StoB_REQ2_p & v87edbb | !StoB_REQ2_p & v872d35;
assign v87ec0b = BtoS_ACK1_p & v879395 | !BtoS_ACK1_p & v87ed0b;
assign v868af8 = BtoS_ACK2_p & v872f79 | !BtoS_ACK2_p & v87e86b;
assign v8730c6 = StoB_REQ2_p & v87ed48 | !StoB_REQ2_p & v85ab45;
assign v87ec46 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v87ee04;
assign v87ecd2 = BtoS_ACK1_p & v8733e9 | !BtoS_ACK1_p & v87ecef;
assign v87ec7a = ENQ_p & v87ec28 | !ENQ_p & v8589e8;
assign v856718 = StoB_REQ0_p & v872e7f | !StoB_REQ0_p & v858bc4;
assign v8731fb = jx0_p & v873741 | !jx0_p & v844f91;
assign v868b41 = BtoS_ACK0_p & v844f99 | !BtoS_ACK0_p & v872fb2;
assign v872b5c = BtoS_ACK0_p & v87ed62 | !BtoS_ACK0_p & v872e9a;
assign BtoS_ACK1_n = !v87df27;
assign v87ec35 = BtoS_ACK0_p & v87edd1 | !BtoS_ACK0_p & v8731cf;
assign v87ed9f = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & v87edcb;
assign v87ed3b = StoB_REQ2_p & v868aba | !StoB_REQ2_p & v87286f;
assign v8598e6 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v87ebe4;
assign jx2_n = v872b76;
assign v858f67 = stateG7_0_p & v8733de | !stateG7_0_p & v87ec89;
assign v87ec1d = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v8728b4;
assign v874242 = BtoS_ACK3_p & v857ea2 | !BtoS_ACK3_p & v8733e9;
assign v868b0e = DEQ_p & v8732f1 | !DEQ_p & v872de2;
assign v87eceb = BtoS_ACK2_p & v87ec96 | !BtoS_ACK2_p & v8731d4;
assign v872837 = BtoS_ACK2_p & v87ecbb | !BtoS_ACK2_p & v8750ad;
assign v87ecb6 = EMPTY_p & v868b6d | !EMPTY_p & v868adc;
assign v8737a3 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v87ef9b;
assign v876238 = stateG12_p & v873307 | !stateG12_p & v872ec6;
assign v872927 = BtoS_ACK2_p & v872f67 | !BtoS_ACK2_p & v8737c6;
assign v87e86b = StoB_REQ2_p & v87eeaa | !StoB_REQ2_p & v873379;
assign v852eb2 = BtoS_ACK1_p & v87ed62 | !BtoS_ACK1_p & v87ed80;
assign v87378d = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87ebee;
assign v8728c0 = DEQ_p & v87ec95 | !DEQ_p & v87edb3;
assign v8732c2 = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v87ec71;
assign v87ed01 = jx0_p & v874c37 | !jx0_p & v844f91;
assign v87459e = DEQ_p & v872f1f | !DEQ_p & v873126;
assign v858aae = StoB_REQ1_p & v844fa9 | !StoB_REQ1_p & v873071;
assign v87ece6 = FULL_p & v87eca9 | !FULL_p & v872d50;
assign v873079 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v85448e;
assign v87ec56 = StoB_REQ1_p & v868aba | !StoB_REQ1_p & v87ed6b;
assign v872cd4 = EMPTY_p & v872b6a | !EMPTY_p & !v844f91;
assign v854114 = BtoS_ACK0_p & v8727fb | !BtoS_ACK0_p & v8736d4;
assign v87ec0a = StoB_REQ1_p & v87ed2f | !StoB_REQ1_p & v87ed3f;
assign v87ec97 = DEQ_p & v872c73 | !DEQ_p & v85884d;
assign v8567f5 = BtoS_ACK0_p & v87ed1e | !BtoS_ACK0_p & v872dbf;
assign v85409b = stateG7_1_p & v844f9f | !stateG7_1_p & v844f91;
assign jx1_n = !v87aed9;
assign v87322c = BtoS_ACK2_p & v859541 | !BtoS_ACK2_p & v855989;
assign v87ec3d = jx1_p & v87ef7a | !jx1_p & v85259e;
assign v8757d4 = EMPTY_p & v87eccc | !EMPTY_p & v872878;
assign v8538fd = StoB_REQ3_p & v868aba | !StoB_REQ3_p & v844f91;
assign v87377f = ENQ_p & v868b92 | !ENQ_p & v873774;
assign v87ed97 = BtoS_ACK2_p & v858d4f | !BtoS_ACK2_p & v868b3d;
assign v872f69 = StoB_REQ2_p & v872de4 | !StoB_REQ2_p & v87ecd7;
assign v875270 = BtoS_ACK1_p & v868aba | !BtoS_ACK1_p & v87ec55;
assign v852e67 = stateG7_1_p & v844f91 | !stateG7_1_p & v844f9f;
assign v8733ec = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & !v87eef6;
assign v872d35 = StoB_REQ3_p & v87338a | !StoB_REQ3_p & !v868aba;
assign v87ec60 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v873383;
assign v87e8f4 = jx1_p & v874c36 | !jx1_p & v87459e;
assign v872c17 = BtoS_ACK0_p & v87ed83 | !BtoS_ACK0_p & v872fee;
assign v85724c = StoB_REQ0_p & v872c51 | !StoB_REQ0_p & v87ec48;
assign v87ee04 = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & !v844f9b;
assign v872c10 = BtoS_ACK1_p & v873375 | !BtoS_ACK1_p & v8728da;
assign v8745a5 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v87ec2c;
assign v857022 = BtoS_ACK0_p & v87ef9b | !BtoS_ACK0_p & v87edd3;
assign v853e70 = DEQ_p & v852613 | !DEQ_p & v844fa5;
assign v873238 = BtoS_ACK0_p & v872f14 | !BtoS_ACK0_p & v858cf2;
assign v87ecbb = StoB_REQ2_p & v8750ad | !StoB_REQ2_p & v844f91;
assign v875285 = EMPTY_p & v87ed71 | !EMPTY_p & v844f91;
assign v855c35 = BtoS_ACK0_p & v87ec1a | !BtoS_ACK0_p & v87ed7b;
assign v872de2 = EMPTY_p & v874047 | !EMPTY_p & v8732f1;
assign v87ecc6 = BtoS_ACK1_p & v872c60 | !BtoS_ACK1_p & v87ed80;
assign v872ee2 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v859947;
assign v87e8ce = BtoS_ACK0_p & v8728da | !BtoS_ACK0_p & v87eee5;
assign v872fbc = StoB_REQ2_p & v872c60 | !StoB_REQ2_p & v844f91;
assign v872835 = DEQ_p & v844f91 | !DEQ_p & v872d64;
assign v868af3 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & v8752b0;
assign v872fc4 = BtoS_ACK0_p & v87eca5 | !BtoS_ACK0_p & v8730d5;
assign v859a0a = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v873227;
assign v873169 = EMPTY_p & v872d50 | !EMPTY_p & v844f91;
assign v87ed79 = stateG7_0_p & v844f91 | !stateG7_0_p & v852e67;
assign v87e8df = BtoS_ACK2_p & v856f49 | !BtoS_ACK2_p & v87e855;
assign v87ef9a = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844f97;
assign v872f42 = FULL_p & v87ecb2 | !FULL_p & v872f1f;
assign v87edb3 = jx0_p & v87ec42 | !jx0_p & v86284b;
assign v874047 = jx0_p & v87ed98 | !jx0_p & !v868b41;
assign v8685f8 = jx1_p & v872ea3 | !jx1_p & !v872c18;
assign v872d56 = BtoS_ACK0_p & v844f9b | !BtoS_ACK0_p & v87ec99;
assign v872822 = EMPTY_p & v872ddf | !EMPTY_p & v844f91;
assign v87e848 = jx1_p & v87edb2 | !jx1_p & v873774;
assign v87ebf3 = jx0_p & v844f9b | !jx0_p & !v87ed71;
assign v844fab = BtoS_ACK3_p & v844f91 | !BtoS_ACK3_p & !v844f91;
assign v873319 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v87332c;
assign v8572b7 = EMPTY_p & v872f47 | !EMPTY_p & v868ae0;
assign v868ac6 = BtoS_ACK0_p & v872f59 | !BtoS_ACK0_p & v87304f;
assign v8731ae = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & v87ec5c;
assign v87ed40 = EMPTY_p & v855c5b | !EMPTY_p & v87ed04;
assign v868bef = jx2_p & v87ec7a | !jx2_p & v872e8e;
assign v87ef71 = EMPTY_p & v872915 | !EMPTY_p & v87ecb3;
assign v862858 = jx2_p & v874051 | !jx2_p & v87ebe9;
assign v87ec70 = BtoS_ACK0_p & v872863 | !BtoS_ACK0_p & v85b0b9;
assign v87edc4 = StoB_REQ2_p & v872d64 | !StoB_REQ2_p & v844f91;
assign v872819 = BtoS_ACK1_p & v87ed5b | !BtoS_ACK1_p & v87ed1c;
assign v873726 = StoB_REQ3_p & v87ec98 | !StoB_REQ3_p & v874242;
assign v875111 = RtoB_ACK0_n & v844f9f | !RtoB_ACK0_n & v85271e;
assign v872d6b = StoB_REQ0_p & v872e81 | !StoB_REQ0_p & v8752b0;
assign v87efcf = BtoS_ACK1_p & v8757ca | !BtoS_ACK1_p & v87ecb5;
assign v872ec6 = BtoS_ACK0_p & v8732c4 | !BtoS_ACK0_p & v8727f7;
assign v872f13 = BtoS_ACK0_p & v87ecea | !BtoS_ACK0_p & v872d64;
assign v868b4a = FULL_p & v87e8d0 | !FULL_p & v87291f;
assign jx0_n = !v87b3e9;
assign v87ec48 = BtoS_ACK1_p & v87eec0 | !BtoS_ACK1_p & v8737ab;
assign v8525dc = DEQ_p & v868b9a | !DEQ_p & v87ecb6;
assign v858363 = StoB_REQ0_p & v85ac62 | !StoB_REQ0_p & v87eda8;
assign v87b3e9 = jx2_p & v844f91 | !jx2_p & !v874063;
assign v852227 = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v872e81;
assign v87ebe9 = ENQ_p & v872df4 | !ENQ_p & v8750bd;
assign v87ed92 = BtoS_ACK2_p & v87ec2d | !BtoS_ACK2_p & v87ed62;
assign v844f95 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & !v844f91;
assign v87ec67 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v87edbb;
assign v872f47 = jx0_p & v87e82a | !jx0_p & v8731b9;
assign v85a741 = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v876307;
assign v872863 = StoB_REQ1_p & v87ed9f | !StoB_REQ1_p & v844f91;
assign v868b29 = StoB_REQ1_p & v8750ad | !StoB_REQ1_p & v8733da;
assign v87e85d = BtoS_ACK1_p & v872c60 | !BtoS_ACK1_p & v872c81;
assign v87eda1 = ENQ_p & v87ef46 | !ENQ_p & v87ec20;
assign v87ef7a = DEQ_p & v87292f | !DEQ_p & v873042;
assign v87ec01 = stateG12_p & v872ff7 | !stateG12_p & v87efcc;
assign v85a712 = BtoS_ACK1_p & v872fa7 | !BtoS_ACK1_p & v85a741;
assign v873723 = StoB_REQ3_p & v87338a | !StoB_REQ3_p & v8757c6;
assign v8588f4 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & v872e81;
assign v852af2 = StoB_REQ2_p & v87338a | !StoB_REQ2_p & !v87ef04;
assign v852d87 = StoB_REQ3_p & v872e81 | !StoB_REQ3_p & v8733e9;
assign v872e80 = BtoS_ACK0_p & v872e99 | !BtoS_ACK0_p & v868b71;
assign v868ba1 = StoB_REQ3_p & v87338a | !StoB_REQ3_p & v874242;
assign v87eeef = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & v844fa9;
assign v8730eb = StoB_REQ1_p & v8750ad | !StoB_REQ1_p & v872837;
assign v87edf9 = StoB_REQ1_p & v86e02d | !StoB_REQ1_p & v844f9d;
assign v87ec82 = StoB_REQ0_p & v872d64 | !StoB_REQ0_p & v844f91;
assign v868aba = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v87eeaa;
assign v873307 = BtoS_ACK0_p & v87ec5a | !BtoS_ACK0_p & v856719;
assign v87ec1c = StoB_REQ3_p & v87ec98 | !StoB_REQ3_p & v8733e9;
assign v872d03 = BtoS_ACK2_p & v87ebe3 | !BtoS_ACK2_p & v8730f3;
assign v852d67 = FULL_p & v873074 | !FULL_p & v868b3a;
assign v87ed47 = StoB_REQ1_p & v87eda9 | !StoB_REQ1_p & v873077;
assign v87ec71 = BtoS_ACK2_p & v872916 | !BtoS_ACK2_p & v857beb;
assign v874df5 = RtoB_ACK0_n & v844f91 | !RtoB_ACK0_n & v87efc2;
assign v8730b0 = BtoS_ACK1_p & v872f69 | !BtoS_ACK1_p & v87ed47;
assign v872916 = StoB_REQ2_p & v872d35 | !StoB_REQ2_p & !v868aba;
assign v873342 = StoB_REQ1_p & v87939c | !StoB_REQ1_p & v872f22;
assign v854111 = StoB_REQ2_p & v8745a5 | !StoB_REQ2_p & v8733e9;
assign v87edbf = jx0_p & v874056 | !jx0_p & v87ed6d;
assign v87eda6 = StoB_REQ2_p & v856f49 | !StoB_REQ2_p & v8745a5;
assign v87ec14 = BtoS_ACK0_p & v87ed62 | !BtoS_ACK0_p & v87ebf4;
assign v876314 = BtoR_REQ1_p & v844f91 | !BtoR_REQ1_p & v844f9f;
assign v87ec98 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & v858f67;
assign v87ece0 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v872830;
assign v87291a = stateG7_0_p & v844f9f | !stateG7_0_p & v85409b;
assign v87ef41 = StoB_REQ0_p & v868b76 | !StoB_REQ0_p & !v872c10;
assign v87ecd5 = EMPTY_p & v87eda4 | !EMPTY_p & v844f91;
assign v87edb0 = jx1_p & v873189 | !jx1_p & !v8732cb;
assign v87ed2d = BtoS_ACK1_p & v87bbdd | !BtoS_ACK1_p & v87622b;
assign v868b8b = StoB_REQ3_p & v856f49 | !StoB_REQ3_p & v8733e9;
assign v874d66 = BtoS_ACK1_p & v87ed55 | !BtoS_ACK1_p & v873342;
assign v87ecfe = DEQ_p & v87ed71 | !DEQ_p & v875285;
assign v8733c1 = StoB_REQ1_p & v859412 | !StoB_REQ1_p & v872db6;
assign v8757ca = StoB_REQ2_p & v87302a | !StoB_REQ2_p & v85ab45;
assign v87edc6 = jx0_p & v872e0f | !jx0_p & v858b3f;
assign v872f5d = StoB_REQ0_p & v872819 | !StoB_REQ0_p & v87372a;
assign v873298 = FULL_p & v87e83a | !FULL_p & v854114;
assign v87ed80 = BtoS_ACK2_p & v87ed62 | !BtoS_ACK2_p & v87eda9;
assign v8728aa = BtoS_ACK1_p & v87eeaa | !BtoS_ACK1_p & v868af8;
assign v872e09 = jx0_p & v872e80 | !jx0_p & v852d93;
assign v872e81 = RtoB_ACK0_p & v844f91 | !RtoB_ACK0_p & !v874df5;
assign v87304f = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v855880;
assign v874226 = jx0_p & v873238 | !jx0_p & v87e7e0;
assign v852626 = StoB_REQ1_p & v87ec2d | !StoB_REQ1_p & v872c81;
assign v87291d = BtoS_ACK0_p & v87ec65 | !BtoS_ACK0_p & v868b13;
assign v87ed13 = StoB_REQ2_p & v8728cb | !StoB_REQ2_p & v87ed27;
assign v873333 = BtoS_ACK2_p & v8737e4 | !BtoS_ACK2_p & v8564be;
assign v87372e = ENQ_p & v872dd8 | !ENQ_p & v87e848;
assign v872dbf = StoB_REQ0_p & v87ecc6 | !StoB_REQ0_p & v87edd7;
assign v87ec3a = EMPTY_p & v87ec04 | !EMPTY_p & !v87edbf;
assign v87ed1e = StoB_REQ1_p & v872c60 | !StoB_REQ1_p & v87ec12;
assign v8733de = stateG7_1_p & v844faf | !stateG7_1_p & v87283c;
assign v872eae = StoB_REQ0_p & v873759 | !StoB_REQ0_p & v87ec0b;
assign v8732c4 = StoB_REQ1_p & v872e81 | !StoB_REQ1_p & v872fa7;
assign v876307 = BtoS_ACK2_p & v873327 | !BtoS_ACK2_p & v87ec05;
assign v87281e = jx0_p & v872f1f | !jx0_p & v872f42;
assign v868aef = BtoS_ACK0_p & v87ec46 | !BtoS_ACK0_p & v87ece0;
assign v873177 = StoB_REQ0_p & v87ebf1 | !StoB_REQ0_p & v87e85b;
assign v872dca = StoB_REQ0_p & v87ee95 | !StoB_REQ0_p & v87efcf;
assign v844f9b = StoB_REQ3_p & v844f91 | !StoB_REQ3_p & !v844f91;
assign v87ed48 = StoB_REQ3_p & v87302a | !StoB_REQ3_p & v87ec98;
assign v8736f8 = BtoS_ACK1_p & v87bbdd | !BtoS_ACK1_p & v87ec56;
assign v873074 = BtoS_ACK0_p & v87ecc3 | !BtoS_ACK0_p & v8793a7;
assign v872d34 = StoB_REQ0_p & v868be9 | !StoB_REQ0_p & v874d66;
assign v8757c6 = BtoS_ACK3_p & v87302a | !BtoS_ACK3_p & v872e81;
assign v87332c = StoB_REQ0_p & v87ec34 | !StoB_REQ0_p & !v844f91;
assign v872f89 = ENQ_p & v87e8f4 | !ENQ_p & !v87ec50;
assign v873172 = StoB_REQ3_p & v872d64 | !StoB_REQ3_p & v844f91;
assign v87eddd = BtoS_ACK2_p & v872fa7 | !BtoS_ACK2_p & v87ec05;
assign v87ee0f = StoB_REQ0_p & v872c60 | !StoB_REQ0_p & v858bae;
assign v872e78 = BtoS_ACK0_p & v87370d | !BtoS_ACK0_p & v872eae;
assign v8598ae = jx1_p & v8737c4 | !jx1_p & v868bac;
assign v87ec08 = StoB_REQ3_p & v87ed9f | !StoB_REQ3_p & v844f91;
assign v868b9a = jx0_p & v8731a1 | !jx0_p & v8567f5;
assign v8757d7 = BtoS_ACK0_p & v8732c4 | !BtoS_ACK0_p & v872d6b;
assign v873779 = BtoS_ACK1_p & v873375 | !BtoS_ACK1_p & v8732c2;
assign v852cab = FULL_p & v87e816 | !FULL_p & v87e83a;
assign v87ed2f = BtoS_ACK2_p & v872e81 | !BtoS_ACK2_p & v8588f4;
assign v87ec1b = StoB_REQ2_p & v844f91 | !StoB_REQ2_p & v872d64;
assign v87ec2a = BtoS_ACK1_p & v87e86b | !BtoS_ACK1_p & v868bde;
assign v87edae = BtoS_ACK0_p & v844f97 | !BtoS_ACK0_p & v87ef9a;
assign v872f14 = StoB_REQ1_p & v868aba | !StoB_REQ1_p & v8728f3;
assign v868b6d = jx0_p & v87ed10 | !jx0_p & v872e78;
assign v87ecb3 = jx0_p & v844f91 | !jx0_p & v87ece6;
assign v87ed45 = StoB_REQ2_p & v857ea2 | !StoB_REQ2_p & v87ed27;
assign v859541 = StoB_REQ2_p & v873723 | !StoB_REQ2_p & v87ec5e;
assign v872949 = StoB_REQ2_p & v872c60 | !StoB_REQ2_p & v87ee84;
assign v87ed15 = jx1_p & v87ec97 | !jx1_p & v87293b;
assign v87ed27 = StoB_REQ3_p & v8733e9 | !StoB_REQ3_p & v844f91;
assign v87ee95 = BtoS_ACK1_p & v87302a | !BtoS_ACK1_p & v872e22;
assign v87ebe3 = StoB_REQ2_p & v87302a | !StoB_REQ2_p & v87ec98;
assign v8736d4 = StoB_REQ0_p & v87338a | !StoB_REQ0_p & !v87df12;
assign v87ec72 = BtoS_ACK0_p & v87ed1e | !BtoS_ACK0_p & v87ee0f;
assign v87370d = StoB_REQ1_p & v857ea2 | !StoB_REQ1_p & v87ee9d;
assign v87eca7 = BtoS_ACK1_p & v844f91 | !BtoS_ACK1_p & !v873071;
assign v868b3a = BtoS_ACK0_p & v872f4c | !BtoS_ACK0_p & v872dca;
assign v8793ad = jx2_p & v876227 | !jx2_p & v87ee8e;
assign v872fb8 = stateG7_0_p & v852e67 | !stateG7_0_p & v85409b;
assign v87df12 = BtoS_ACK1_p & v87edb8 | !BtoS_ACK1_p & !v85a55b;
assign v87ed9d = StoB_REQ1_p & v872e6f | !StoB_REQ1_p & v872d7f;
assign v87ef46 = BtoS_ACK0_p & v844f91 | !BtoS_ACK0_p & !v844fa7;
assign v87e82a = BtoS_ACK0_p & v87ec25 | !BtoS_ACK0_p & v87e8be;
assign v872da9 = StoB_REQ0_p & v844f91 | !StoB_REQ0_p & v87ede2;
assign v872eb0 = BtoS_ACK1_p & v87ec41 | !BtoS_ACK1_p & v87ec15;
assign v844f97 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & !v844f91;
assign v87edd1 = StoB_REQ1_p & v844f91 | !StoB_REQ1_p & v844f99;
assign v872dff = BtoS_ACK2_p & v87302a | !BtoS_ACK2_p & v87edd0;
assign v87ee8e = ENQ_p & v844fa5 | !ENQ_p & !v87ec3d;
assign v8737d6 = jx0_p & v844f9b | !jx0_p & !v868aef;
assign v87ec22 = EMPTY_p & v87ef70 | !EMPTY_p & !v87ec63;
assign v87ee8b = StoB_REQ3_p & v856f49 | !StoB_REQ3_p & v87ecbd;
assign v872f4e = stateG7_1_p & v844faf | !stateG7_1_p & !v844f91;
assign v872fa7 = StoB_REQ2_p & v872e81 | !StoB_REQ2_p & v852d87;
assign v852d6f = StoB_REQ2_p & v87ed5b | !StoB_REQ2_p & v87ec5e;
assign v87ed2c = StoB_REQ3_p & v87eeaa | !StoB_REQ3_p & v87ed6c;
assign v87ed81 = BtoS_ACK1_p & v87bbdd | !BtoS_ACK1_p & v873181;
assign v87ed51 = BtoS_ACK2_p & v872949 | !BtoS_ACK2_p & v872fbc;
assign v87ecbe = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v852af2;
assign v86283e = BtoS_ACK0_p & v8732c4 | !BtoS_ACK0_p & v8757c5;
assign v87ed76 = StoB_REQ2_p & v87ef9c | !StoB_REQ2_p & v872ed3;
assign v85260c = StoB_REQ1_p & v87ed80 | !StoB_REQ1_p & v872f69;
assign v872830 = BtoS_ACK1_p & v844f99 | !BtoS_ACK1_p & v87ec46;
assign v874051 = ENQ_p & v872835 | !ENQ_p & v8750bd;
assign v872c93 = StoB_REQ0_p & v852eb2 | !StoB_REQ0_p & v873048;
assign v87ef83 = BtoS_ACK1_p & v87ec41 | !BtoS_ACK1_p & v872927;
assign v87ec15 = StoB_REQ1_p & v87e8df | !StoB_REQ1_p & v87287b;
assign v87ef15 = BtoS_ACK1_p & v868aba | !BtoS_ACK1_p & v87ed68;
assign v858d4f = StoB_REQ2_p & v8564be | !StoB_REQ2_p & v87ec1c;
assign v872f79 = StoB_REQ2_p & v87eeaa | !StoB_REQ2_p & v868aba;
assign v855cab = stateG7_1_p & v873370 | !stateG7_1_p & v844f9f;
assign v876227 = ENQ_p & v853e70 | !ENQ_p & !v87332a;
assign v8731b9 = BtoS_ACK0_p & v87ecdb | !BtoS_ACK0_p & v872fe0;
assign v87ebf1 = BtoS_ACK1_p & v85a673 | !BtoS_ACK1_p & v873333;
assign v87ec99 = BtoS_ACK1_p & v844f9b | !BtoS_ACK1_p & !v844f91;
assign v87ecde = ENQ_p & v87330a | !ENQ_p & v87ed36;
assign v8728da = StoB_REQ1_p & v87338a | !StoB_REQ1_p & v873375;
assign v858b3f = BtoS_ACK0_p & v872d64 | !BtoS_ACK0_p & v87eee0;
assign v87ec5e = StoB_REQ3_p & v87338a | !StoB_REQ3_p & v8733e9;
assign v872c73 = jx0_p & v87291d | !jx0_p & v8598fe;
assign v879392 = DEQ_p & v844fb9 | !DEQ_p & !v87eee6;
assign v8732c5 = StoB_REQ2_p & v868ace | !StoB_REQ2_p & v8538fd;
assign v872d0b = BtoS_ACK0_p & v873375 | !BtoS_ACK0_p & v87ec8e;
assign v8594bd = DEQ_p & v872e09 | !DEQ_p & v8572b7;
assign v868bac = jx0_p & v857e91 | !jx0_p & !v844f91;
assign v872e92 = StoB_REQ0_p & v87ec2d | !StoB_REQ0_p & v872e9a;
assign v87ed1c = BtoS_ACK2_p & v872e8b | !BtoS_ACK2_p & v873723;
assign v872ed3 = StoB_REQ3_p & v857ea2 | !StoB_REQ3_p & v844f91;
assign v872f60 = stateG12_p & v873307 | !stateG12_p & v86283e;
assign v872d64 = RtoB_ACK0_p & v844fad | !RtoB_ACK0_p & v87283c;
assign v87332b = BtoS_ACK1_p & v87ec12 | !BtoS_ACK1_p & v85260c;
assign SLC0_n = (jx0_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))) | (!jx0_n & ((jx1_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))) | (!jx1_n & ((jx2_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))) | (!jx2_n & ((EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((StoB_REQ1_n & ((!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))) | (!StoB_REQ1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))) | (!StoB_REQ0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n)))))))))))))))))))))))));
assign ENQ_n = (EMPTY_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))))) | (!stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n & ((!DEQ_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!DEQ_n))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n & ((DEQ_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((DEQ_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((DEQ_n))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))))))))))))))) | (!FULL_n & ((stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n))) | (!BtoS_ACK1_n & ((SLC0_n) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n))))))))))) | (!stateG12_n & ((BtoS_ACK0_n & ((StoB_REQ0_n & ((!DEQ_n))))) | (!BtoS_ACK0_n & ((BtoS_ACK1_n & ((StoB_REQ1_n & ((!DEQ_n))))) | (!BtoS_ACK1_n & ((SLC0_n & ((!DEQ_n))) | (!SLC0_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n)))))))))))))))));
assign SLC1_n = (jx0_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))))) | (!jx0_n & ((jx1_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))))) | (!jx1_n & ((jx2_n & ((EMPTY_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))))) | (!jx2_n & ((EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))))))) | (!EMPTY_n & ((FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))) | (!StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((DEQ_n))))))))))))))))))) | (!FULL_n & ((stateG12_n & ((!BtoS_ACK0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n))))))))))))) | (!stateG12_n & ((!BtoS_ACK0_n & ((StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))) | (!StoB_REQ1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))))))))) | (!StoB_REQ0_n & ((!BtoS_ACK1_n & ((StoB_REQ2_n & ((BtoS_ACK2_n & ((!DEQ_n))) | (!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n))))))))) | (!StoB_REQ2_n & ((!BtoS_ACK2_n & ((BtoS_ACK3_n & ((StoB_REQ3_n & ((!DEQ_n)))))))))))))))))))))))))));
    initial begin
  StoB_REQ0_p = 0;
  StoB_REQ1_p = 0;
  StoB_REQ2_p = 0;
  StoB_REQ3_p = 0;
  RtoB_ACK0_p = 0;
  RtoB_ACK1_p = 0;
  FULL_p = 0;
  EMPTY_p = 1;
  BtoS_ACK0_p = 0;
  BtoS_ACK1_p = 0;
  BtoS_ACK2_p = 0;
  BtoS_ACK3_p = 0;
  BtoR_REQ0_p = 0;
  BtoR_REQ1_p = 0;
  stateG7_0_p = 0;
  stateG7_1_p = 1;
  ENQ_p = 0;
  DEQ_p = 0;
  stateG12_p = 0;
  SLC0_p = 0;
  SLC1_p = 0;
  jx0_p = 0;
  jx1_p = 0;
  jx2_p = 0;
    end
    always @(posedge clock) begin
  StoB_REQ0_p = StoB_REQ0_n;
  StoB_REQ1_p = StoB_REQ1_n;
  StoB_REQ2_p = StoB_REQ2_n;
  StoB_REQ3_p = StoB_REQ3_n;
  RtoB_ACK0_p = RtoB_ACK0_n;
  RtoB_ACK1_p = RtoB_ACK1_n;
  FULL_p = FULL_n;
  EMPTY_p = EMPTY_n;
  BtoS_ACK0_p = BtoS_ACK0_n;
  BtoS_ACK1_p = BtoS_ACK1_n;
  BtoS_ACK2_p = BtoS_ACK2_n;
  BtoS_ACK3_p = BtoS_ACK3_n;
  BtoR_REQ0_p = BtoR_REQ0_n;
  BtoR_REQ1_p = BtoR_REQ1_n;
  stateG7_0_p = stateG7_0_n;
  stateG7_1_p = stateG7_1_n;
  ENQ_p = ENQ_n;
  DEQ_p = DEQ_n;
  stateG12_p = stateG12_n;
  SLC0_p = SLC0_n;
  SLC1_p = SLC1_n;
  jx0_p = jx0_n;
  jx1_p = jx1_n;
  jx2_p = jx2_n;
    end


  DBW7 G7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
  DBW12 G12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
endmodule

//Note that the DBW for G7 works only for two receivers.
module DBW7(stateG7_1_n, stateG7_0_n, stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p);
	input  stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	output stateG7_1_n, stateG7_0_n;
	wire    stateG7_1_p, stateG7_0_p, BtoR_REQ0_p, BtoR_REQ1_p;
	wire    stateG7_1_n, stateG7_0_n;

	assign  stateG7_1_n = (!stateG7_1_p && !BtoR_REQ0_p &&  BtoR_REQ1_p)||
	                      ( stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p)||
	                      ( stateG7_1_p && !stateG7_0_p && !BtoR_REQ0_p && BtoR_REQ1_p);
	assign  stateG7_0_n = (!stateG7_1_p && !BtoR_REQ0_p && !BtoR_REQ1_p);
endmodule
module DBW12(stateG12_n, stateG12_p, EMPTY_p, DEQ_p);
	input  stateG12_p, EMPTY_p, DEQ_p;
	output stateG12_n;
	wire    stateG12_n, stateG12_p, EMPTY_p, DEQ_p;

	assign  stateG12_n = (!stateG12_p && !DEQ_p && !EMPTY_p)||
	                     ( stateG12_p && !DEQ_p);
endmodule
